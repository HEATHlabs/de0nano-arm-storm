-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
--				MEM_SIZE      : natural := 1024;  -- memory cells
--				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				MEM_SIZE      : natural := 2048;  -- memory cells
				LOG2_MEM_SIZE : natural := 11;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
-- bootloader_sdram
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
000000 => x"EA000006",
000001 => x"EAFFFFFE",
000002 => x"EAFFFFFE",
000003 => x"EAFFFFFE",
000004 => x"EAFFFFFE",
000005 => x"E1A00000",
000006 => x"EAFFFFFE",
000007 => x"EAFFFFFE",
000008 => x"E59F0040",
000009 => x"E10F1000",
000010 => x"E3C1107F",
000011 => x"E38110DF",
000012 => x"E129F001",
000013 => x"E1A0D000",
000014 => x"E3A00000",
000015 => x"E1A01000",
000016 => x"E1A02000",
000017 => x"E1A0B000",
000018 => x"E1A07000",
000019 => x"E59FA018",
000020 => x"E1A0E00F",
000021 => x"E1A0F00A",
000022 => x"E1A04000",
000023 => x"E3A00000",
000024 => x"E1A0F004",
000025 => x"EAFFFFFE",
000026 => x"00002000",
000027 => x"000107B0",
000028 => x"E3E03A0F",
000029 => x"E5131FFB",
000030 => x"E20020FF",
000031 => x"E3A00001",
000032 => x"E0010210",
000033 => x"E1A0F00E",
000034 => x"E3E03A0F",
000035 => x"E5130FFB",
000036 => x"E1A0F00E",
000037 => x"E3E01A0F",
000038 => x"E5113FFF",
000039 => x"E20000FF",
000040 => x"E3A02001",
000041 => x"E1833012",
000042 => x"E5013FFF",
000043 => x"E1A0F00E",
000044 => x"E20000FF",
000045 => x"E3A02001",
000046 => x"E1A02012",
000047 => x"E3E01A0F",
000048 => x"E5113FFF",
000049 => x"E1E02002",
000050 => x"E0033002",
000051 => x"E5013FFF",
000052 => x"E1A0F00E",
000053 => x"E3E01A0F",
000054 => x"E5113FFF",
000055 => x"E20000FF",
000056 => x"E3A02001",
000057 => x"E0233012",
000058 => x"E5013FFF",
000059 => x"E1A0F00E",
000060 => x"E3E03A0F",
000061 => x"E5030FFF",
000062 => x"E1A0F00E",
000063 => x"E20000FF",
000064 => x"E3500007",
000065 => x"E92D4010",
000066 => x"E3A0C000",
000067 => x"E3E0E0FF",
000068 => x"E20110FF",
000069 => x"8A000011",
000070 => x"E2403004",
000071 => x"E20330FF",
000072 => x"E3500003",
000073 => x"E1A0E183",
000074 => x"E3E04A0F",
000075 => x"E1A0C180",
000076 => x"9A000007",
000077 => x"E3A030FF",
000078 => x"E1A03E13",
000079 => x"E5142F8B",
000080 => x"E1E03003",
000081 => x"E0022003",
000082 => x"E1822E11",
000083 => x"E5042F8B",
000084 => x"E8BD8010",
000085 => x"E3A030FF",
000086 => x"E1A03C13",
000087 => x"E1E0E003",
000088 => x"E3E02A0F",
000089 => x"E5123F8F",
000090 => x"E003300E",
000091 => x"E1833C11",
000092 => x"E5023F8F",
000093 => x"E8BD8010",
000094 => x"E20000FF",
000095 => x"E3500007",
000096 => x"E3A02000",
000097 => x"8A00000A",
000098 => x"E2403004",
000099 => x"E3500003",
000100 => x"E20320FF",
000101 => x"9A000005",
000102 => x"E3E03A0F",
000103 => x"E5130F8B",
000104 => x"E1A02182",
000105 => x"E1A00230",
000106 => x"E20000FF",
000107 => x"E1A0F00E",
000108 => x"E1A02180",
000109 => x"E3E03A0F",
000110 => x"E5130F8F",
000111 => x"E1A00230",
000112 => x"E20000FF",
000113 => x"E1A0F00E",
000114 => x"E3E02A0F",
000115 => x"E5123FE3",
000116 => x"E3130002",
000117 => x"E3E00000",
000118 => x"15120FE7",
000119 => x"E1A0F00E",
000120 => x"E3E02A0F",
000121 => x"E5123FE3",
000122 => x"E3130001",
000123 => x"0AFFFFFC",
000124 => x"E20030FF",
000125 => x"E5023FE7",
000126 => x"E1A0F00E",
000127 => x"E20000FF",
000128 => x"E3500001",
000129 => x"E3812B01",
000130 => x"03E03A0F",
000131 => x"E3811B09",
000132 => x"13E03A0F",
000133 => x"05031FCF",
000134 => x"15032FCF",
000135 => x"E1A0F00E",
000136 => x"E3E03A0F",
000137 => x"E5030FCB",
000138 => x"E1A0F00E",
000139 => x"E3E02A0F",
000140 => x"E5123FCF",
000141 => x"E3130C01",
000142 => x"1AFFFFFC",
000143 => x"E5020FBF",
000144 => x"E5123FCF",
000145 => x"E3833C01",
000146 => x"E5023FCF",
000147 => x"E3E02A0F",
000148 => x"E5123FCF",
000149 => x"E3130C01",
000150 => x"1AFFFFFC",
000151 => x"E5120FBF",
000152 => x"E1A0F00E",
000153 => x"E3E01A0F",
000154 => x"E5113FC7",
000155 => x"E20000FF",
000156 => x"E3A02001",
000157 => x"E1833012",
000158 => x"E5013FC7",
000159 => x"E1A0F00E",
000160 => x"E20000FF",
000161 => x"E3A02001",
000162 => x"E1A02012",
000163 => x"E3E01A0F",
000164 => x"E5113FC7",
000165 => x"E1E02002",
000166 => x"E0033002",
000167 => x"E5013FC7",
000168 => x"E1A0F00E",
000169 => x"E3E02A0F",
000170 => x"E5123F97",
000171 => x"E1A01420",
000172 => x"E3C33080",
000173 => x"E5023F97",
000174 => x"E5020F9F",
000175 => x"E5021F9B",
000176 => x"E5123F97",
000177 => x"E3833080",
000178 => x"E5023F97",
000179 => x"E1A0F00E",
000180 => x"E92D4030",
000181 => x"E3A0C090",
000182 => x"E20140FE",
000183 => x"E3E0EA0F",
000184 => x"E5DD500F",
000185 => x"E20000FF",
000186 => x"E50E4F93",
000187 => x"E20110FF",
000188 => x"E50ECFAF",
000189 => x"E1A04002",
000190 => x"E203C0FF",
000191 => x"E51E3FAF",
000192 => x"E3130002",
000193 => x"1AFFFFFC",
000194 => x"E51E3FAF",
000195 => x"E3130080",
000196 => x"13E00000",
000197 => x"18BD8030",
000198 => x"E35C0000",
000199 => x"0A000012",
000200 => x"E24C3001",
000201 => x"E203C0FF",
000202 => x"E35C0001",
000203 => x"01A02424",
000204 => x"03E03A0F",
000205 => x"13E03A0F",
000206 => x"05032F93",
000207 => x"15034F93",
000208 => x"E3E02A0F",
000209 => x"E3A03010",
000210 => x"E5023FAF",
000211 => x"E5123FAF",
000212 => x"E3130002",
000213 => x"1AFFFFFC",
000214 => x"E5123FAF",
000215 => x"E3130080",
000216 => x"0AFFFFEC",
000217 => x"E3E00001",
000218 => x"E8BD8030",
000219 => x"E3500077",
000220 => x"1A00000C",
000221 => x"E3E03A0F",
000222 => x"E3A02050",
000223 => x"E5035F93",
000224 => x"E5032FAF",
000225 => x"E1A02003",
000226 => x"E5123FAF",
000227 => x"E3130002",
000228 => x"1AFFFFFC",
000229 => x"E5123FAF",
000230 => x"E2130080",
000231 => x"08BD8030",
000232 => x"E3E00002",
000233 => x"E8BD8030",
000234 => x"E3500072",
000235 => x"13E00003",
000236 => x"18BD8030",
000237 => x"E3813001",
000238 => x"E3E02A0F",
000239 => x"E3A01090",
000240 => x"E5023F93",
000241 => x"E5021FAF",
000242 => x"E5123FAF",
000243 => x"E3130002",
000244 => x"1AFFFFFC",
000245 => x"E5123FAF",
000246 => x"E3130080",
000247 => x"1AFFFFEF",
000248 => x"E3A03068",
000249 => x"E5023FAF",
000250 => x"E3E00A0F",
000251 => x"E5103FAF",
000252 => x"E3130002",
000253 => x"1AFFFFFC",
000254 => x"E5100F93",
000255 => x"E8BD8030",
000256 => x"E20000FF",
000257 => x"E350000F",
000258 => x"979FF100",
000259 => x"EA00000F",
000260 => x"000104D0",
000261 => x"000104C8",
000262 => x"000104C0",
000263 => x"000104B8",
000264 => x"000104B0",
000265 => x"000104A8",
000266 => x"000104A0",
000267 => x"00010498",
000268 => x"00010490",
000269 => x"00010488",
000270 => x"00010480",
000271 => x"00010478",
000272 => x"00010470",
000273 => x"00010468",
000274 => x"00010460",
000275 => x"00010458",
000276 => x"E3A00000",
000277 => x"E1A0F00E",
000278 => x"EE1F0F1F",
000279 => x"E1A0F00E",
000280 => x"EE1E0F1E",
000281 => x"E1A0F00E",
000282 => x"EE1D0F1D",
000283 => x"E1A0F00E",
000284 => x"EE1C0F1C",
000285 => x"E1A0F00E",
000286 => x"EE1B0F1B",
000287 => x"E1A0F00E",
000288 => x"EE1A0F1A",
000289 => x"E1A0F00E",
000290 => x"EE190F19",
000291 => x"E1A0F00E",
000292 => x"EE180F18",
000293 => x"E1A0F00E",
000294 => x"EE170F17",
000295 => x"E1A0F00E",
000296 => x"EE160F16",
000297 => x"E1A0F00E",
000298 => x"EE150F15",
000299 => x"E1A0F00E",
000300 => x"EE140F14",
000301 => x"E1A0F00E",
000302 => x"EE130F13",
000303 => x"E1A0F00E",
000304 => x"EE120F12",
000305 => x"E1A0F00E",
000306 => x"EE110F11",
000307 => x"E1A0F00E",
000308 => x"EE100F10",
000309 => x"E1A0F00E",
000310 => x"E20110FF",
000311 => x"E2411006",
000312 => x"E3510007",
000313 => x"979FF101",
000314 => x"EA000008",
000315 => x"00010514",
000316 => x"00010510",
000317 => x"00010510",
000318 => x"00010510",
000319 => x"00010510",
000320 => x"0001051C",
000321 => x"00010524",
000322 => x"0001050C",
000323 => x"EE0D0F1D",
000324 => x"E1A0F00E",
000325 => x"EE060F16",
000326 => x"E1A0F00E",
000327 => x"EE0B0F1B",
000328 => x"E1A0F00E",
000329 => x"EE0C0F1C",
000330 => x"E1A0F00E",
000331 => x"E92D4010",
000332 => x"E1A04000",
000333 => x"E5D00000",
000334 => x"E3500000",
000335 => x"1A000003",
000336 => x"EA000005",
000337 => x"E5F40001",
000338 => x"E3500000",
000339 => x"0A000002",
000340 => x"EBFFFF22",
000341 => x"E3500000",
000342 => x"CAFFFFF9",
000343 => x"E1A00004",
000344 => x"E8BD8010",
000345 => x"E92D4070",
000346 => x"E2514000",
000347 => x"E1A05000",
000348 => x"E20260FF",
000349 => x"D8BD8070",
000350 => x"EBFFFF12",
000351 => x"E3700001",
000352 => x"E20030FF",
000353 => x"0A000005",
000354 => x"E3560001",
000355 => x"E5C53000",
000356 => x"E1A00003",
000357 => x"E2855001",
000358 => x"0A000003",
000359 => x"E2444001",
000360 => x"E3540000",
000361 => x"CAFFFFF3",
000362 => x"E8BD8070",
000363 => x"EBFFFF0B",
000364 => x"EAFFFFF9",
000365 => x"E92D4030",
000366 => x"E2514000",
000367 => x"E1A05000",
000368 => x"D8BD8030",
000369 => x"E4D50001",
000370 => x"EBFFFF04",
000371 => x"E2544001",
000372 => x"1AFFFFFB",
000373 => x"E8BD8030",
000374 => x"E92D4010",
000375 => x"E20240FF",
000376 => x"E3540008",
000377 => x"83A04008",
000378 => x"8A000001",
000379 => x"E3540000",
000380 => x"03A04001",
000381 => x"E1A02001",
000382 => x"E1A0E004",
000383 => x"E1A0310E",
000384 => x"E35E0001",
000385 => x"E2433004",
000386 => x"E1A0C000",
000387 => x"81A0C330",
000388 => x"E24E3001",
000389 => x"E20CC00F",
000390 => x"E203E0FF",
000391 => x"E35C0009",
000392 => x"E28C3030",
000393 => x"828C3037",
000394 => x"E35E0000",
000395 => x"E4C23001",
000396 => x"1AFFFFF1",
000397 => x"E2443001",
000398 => x"E20330FF",
000399 => x"E0813003",
000400 => x"E5C3E001",
000401 => x"E8BD8010",
000402 => x"E92D4010",
000403 => x"E1A04000",
000404 => x"E3540007",
000405 => x"E3A01010",
000406 => x"E3A00001",
000407 => x"9A000001",
000408 => x"E3A00000",
000409 => x"E8BD8010",
000410 => x"EBFFFEE3",
000411 => x"E3A00006",
000412 => x"EBFFFEFB",
000413 => x"E3A00000",
000414 => x"EBFFFEEB",
000415 => x"E1A00584",
000416 => x"E8BD4010",
000417 => x"EAFFFEE8",
000418 => x"E0603280",
000419 => x"E0800103",
000420 => x"E0800100",
000421 => x"E1A00200",
000422 => x"E3500000",
000423 => x"D1A0F00E",
000424 => x"E1A00000",
000425 => x"E2500001",
000426 => x"1AFFFFFC",
000427 => x"E1A0F00E",
000428 => x"E212C0FF",
000429 => x"0A00000B",
000430 => x"E5D02000",
000431 => x"E5D13000",
000432 => x"E1520003",
000433 => x"0A000004",
000434 => x"EA000008",
000435 => x"E5F02001",
000436 => x"E5F13001",
000437 => x"E1520003",
000438 => x"1A000004",
000439 => x"E24C3001",
000440 => x"E213C0FF",
000441 => x"1AFFFFF8",
000442 => x"E3A00001",
000443 => x"E1A0F00E",
000444 => x"E3A00000",
000445 => x"E1A0F00E",
000446 => x"E92D4030",
000447 => x"E1A04081",
000448 => x"E3540000",
000449 => x"E1A05000",
000450 => x"D3A00000",
000451 => x"D8BD8030",
000452 => x"E3A00000",
000453 => x"E1A01000",
000454 => x"E7D12005",
000455 => x"E2423030",
000456 => x"E082C200",
000457 => x"E3530009",
000458 => x"E242E041",
000459 => x"924C0030",
000460 => x"9A000007",
000461 => x"E0823200",
000462 => x"E35E0005",
000463 => x"E242C061",
000464 => x"92430037",
000465 => x"9A000002",
000466 => x"E0823200",
000467 => x"E35C0005",
000468 => x"92430057",
000469 => x"E2811001",
000470 => x"E1510004",
000471 => x"1AFFFFED",
000472 => x"E8BD8030",
000473 => x"E5D03003",
000474 => x"E5D02002",
000475 => x"E5D01000",
000476 => x"E1833402",
000477 => x"E5D00001",
000478 => x"E1833C01",
000479 => x"E1830800",
000480 => x"E1A0F00E",
000481 => x"E52DE004",
000482 => x"E59F0014",
000483 => x"EBFFFF66",
000484 => x"E59F0010",
000485 => x"EBFFFF64",
000486 => x"E59F000C",
000487 => x"E49DE004",
000488 => x"EAFFFF61",
000489 => x"00011184",
000490 => x"000111E8",
000491 => x"0001124C",
000492 => x"E92D47F0",
000493 => x"E3A00000",
000494 => x"E24DD014",
000495 => x"EBFFFE4B",
000496 => x"E3A0100D",
000497 => x"E3A000C3",
000498 => x"EBFFFF42",
000499 => x"E3A00063",
000500 => x"EBFFFEB3",
000501 => x"E3A00006",
000502 => x"EBFFFF08",
000503 => x"E3A01006",
000504 => x"E3C00008",
000505 => x"EBFFFF3B",
000506 => x"E3A0000D",
000507 => x"EBFFFF03",
000508 => x"E1A008A0",
000509 => x"E1E00000",
000510 => x"E200000F",
000511 => x"E3500001",
000512 => x"03A04030",
000513 => x"028DA006",
000514 => x"028D900F",
000515 => x"0A000020",
000516 => x"E3500002",
000517 => x"0A00007E",
000518 => x"E59F085C",
000519 => x"EBFFFF42",
000520 => x"E59F0858",
000521 => x"EBFFFF40",
000522 => x"E59F0854",
000523 => x"EBFFFF3E",
000524 => x"E59F0850",
000525 => x"EBFFFF3C",
000526 => x"E59F084C",
000527 => x"EBFFFF3A",
000528 => x"E59F0848",
000529 => x"EBFFFF38",
000530 => x"E59F0844",
000531 => x"EBFFFF36",
000532 => x"E59F0840",
000533 => x"EBFFFF34",
000534 => x"E28DA006",
000535 => x"E59F0838",
000536 => x"EBFFFF31",
000537 => x"E1A0100A",
000538 => x"E3A02008",
000539 => x"E3A00401",
000540 => x"EBFFFF58",
000541 => x"E1A0000A",
000542 => x"EBFFFF2B",
000543 => x"E59F081C",
000544 => x"EBFFFF29",
000545 => x"EBFFFFBE",
000546 => x"E28D900F",
000547 => x"EBFFFE4D",
000548 => x"E1A04000",
000549 => x"E3A0000D",
000550 => x"EBFFFED8",
000551 => x"E3100801",
000552 => x"03A06001",
000553 => x"03A050A0",
000554 => x"1A00003D",
000555 => x"E3A04000",
000556 => x"E59F07EC",
000557 => x"EBFFFF1C",
000558 => x"E1A01005",
000559 => x"E1A02004",
000560 => x"E3A03002",
000561 => x"E3A00072",
000562 => x"E58D4000",
000563 => x"EBFFFE7F",
000564 => x"E1A01005",
000565 => x"E5CD000F",
000566 => x"E3A02001",
000567 => x"E3A03002",
000568 => x"E3A00072",
000569 => x"E58D4000",
000570 => x"EBFFFE78",
000571 => x"E3A02002",
000572 => x"E1A03002",
000573 => x"E5CD0010",
000574 => x"E1A01005",
000575 => x"E3A00072",
000576 => x"E58D4000",
000577 => x"EBFFFE71",
000578 => x"E3A03002",
000579 => x"E5CD0011",
000580 => x"E1A01005",
000581 => x"E3A00072",
000582 => x"E3A02003",
000583 => x"E58D4000",
000584 => x"EBFFFE6A",
000585 => x"E5DD300F",
000586 => x"E20000FF",
000587 => x"E3530053",
000588 => x"E5CD0012",
000589 => x"1A000002",
000590 => x"E5DD3010",
000591 => x"E353004D",
000592 => x"0A00006B",
000593 => x"E59F075C",
000594 => x"EBFFFEF7",
000595 => x"E3560000",
000596 => x"0AFFFFCD",
000597 => x"E59F0750",
000598 => x"EBFFFEF3",
000599 => x"E3A0100D",
000600 => x"E3A00000",
000601 => x"EBFFFEDB",
000602 => x"E3A00006",
000603 => x"EBFFFEA3",
000604 => x"E3A01006",
000605 => x"E3C00008",
000606 => x"EBFFFED6",
000607 => x"E3A00006",
000608 => x"EBFFFE9E",
000609 => x"E1E00000",
000610 => x"E2000002",
000611 => x"E1E00000",
000612 => x"E3A01006",
000613 => x"EBFFFECF",
000614 => x"E3A00401",
000615 => x"EBFFFDAD",
000616 => x"EAFFFFFE",
000617 => x"E3540034",
000618 => x"0A000029",
000619 => x"CA00001C",
000620 => x"E3540031",
000621 => x"0A000036",
000622 => x"DA000098",
000623 => x"E3540032",
000624 => x"0A0000A2",
000625 => x"E3540033",
000626 => x"1A000098",
000627 => x"E1A00004",
000628 => x"EBFFFE02",
000629 => x"E59F06D4",
000630 => x"EBFFFED3",
000631 => x"E1A00009",
000632 => x"E3A01002",
000633 => x"E3A02001",
000634 => x"EBFFFEDD",
000635 => x"E3A01002",
000636 => x"E1A00009",
000637 => x"EBFFFF3F",
000638 => x"E21010FF",
000639 => x"11A05001",
000640 => x"13A06000",
000641 => x"1AFFFFA8",
000642 => x"E59F06A4",
000643 => x"EBFFFEC6",
000644 => x"EAFFFF9D",
000645 => x"E3A04033",
000646 => x"E28DA006",
000647 => x"E28D900F",
000648 => x"EAFFFF9B",
000649 => x"E3540066",
000650 => x"0A00002A",
000651 => x"DA0000AD",
000652 => x"E3540068",
000653 => x"0A00010F",
000654 => x"E3540072",
000655 => x"1A00007B",
000656 => x"E1A00004",
000657 => x"EBFFFDE5",
000658 => x"E3A006FF",
000659 => x"E280F20F",
000660 => x"EAFFFFFE",
000661 => x"E1A00004",
000662 => x"EBFFFDE0",
000663 => x"E59F064C",
000664 => x"EBFFFEB1",
000665 => x"E1A00009",
000666 => x"E3A01002",
000667 => x"E3A02001",
000668 => x"EBFFFEBB",
000669 => x"E1A00009",
000670 => x"E3A01002",
000671 => x"EBFFFF1D",
000672 => x"E21080FF",
000673 => x"1A0000A4",
000674 => x"E59F0628",
000675 => x"EBFFFEA6",
000676 => x"EAFFFF7D",
000677 => x"E1A00004",
000678 => x"EBFFFDD0",
000679 => x"E59F0618",
000680 => x"EBFFFEA1",
000681 => x"E1A00009",
000682 => x"E3A01004",
000683 => x"E3A02000",
000684 => x"EBFFFEAB",
000685 => x"E5DD300F",
000686 => x"E3530053",
000687 => x"1A000002",
000688 => x"E5DD3010",
000689 => x"E353004D",
000690 => x"0A000115",
000691 => x"E59F05EC",
000692 => x"EBFFFE95",
000693 => x"EAFFFF6C",
000694 => x"E1A00004",
000695 => x"EBFFFDBF",
000696 => x"E59F05DC",
000697 => x"EBFFFE90",
000698 => x"E59F05D8",
000699 => x"EBFFFE8E",
000700 => x"EAFFFF65",
000701 => x"E5DD3011",
000702 => x"E3530042",
000703 => x"1AFFFF90",
000704 => x"E3500052",
000705 => x"1AFFFF8E",
000706 => x"E1A01005",
000707 => x"E3A02004",
000708 => x"E2433040",
000709 => x"E2800020",
000710 => x"E58D4000",
000711 => x"EBFFFDEB",
000712 => x"E1A01005",
000713 => x"E5CD000F",
000714 => x"E3A02005",
000715 => x"E3A03002",
000716 => x"E3A00072",
000717 => x"E58D4000",
000718 => x"EBFFFDE4",
000719 => x"E1A01005",
000720 => x"E5CD0010",
000721 => x"E3A02006",
000722 => x"E3A03002",
000723 => x"E3A00072",
000724 => x"E58D4000",
000725 => x"EBFFFDDD",
000726 => x"E1A01005",
000727 => x"E5CD0011",
000728 => x"E3A02007",
000729 => x"E3A03002",
000730 => x"E3A00072",
000731 => x"E58D4000",
000732 => x"EBFFFDD6",
000733 => x"E5CD0012",
000734 => x"E1A00009",
000735 => x"EBFFFEF8",
000736 => x"E2907004",
000737 => x"0A000022",
000738 => x"E1A06004",
000739 => x"E2842008",
000740 => x"E1A01005",
000741 => x"E3A03002",
000742 => x"E3A00072",
000743 => x"E58D6000",
000744 => x"EBFFFDCA",
000745 => x"E2842009",
000746 => x"E5CD000F",
000747 => x"E1A01005",
000748 => x"E3A03002",
000749 => x"E3A00072",
000750 => x"E58D6000",
000751 => x"EBFFFDC3",
000752 => x"E284200A",
000753 => x"E5CD0010",
000754 => x"E1A01005",
000755 => x"E3A03002",
000756 => x"E3A00072",
000757 => x"E58D6000",
000758 => x"EBFFFDBC",
000759 => x"E284200B",
000760 => x"E5CD0011",
000761 => x"E1A01005",
000762 => x"E3A03002",
000763 => x"E3A00072",
000764 => x"E58D6000",
000765 => x"EBFFFDB5",
000766 => x"E5CD0012",
000767 => x"E1A00009",
000768 => x"EBFFFED7",
000769 => x"E4840004",
000770 => x"E1540007",
000771 => x"13540902",
000772 => x"3AFFFFDD",
000773 => x"E59F04B0",
000774 => x"EBFFFE43",
000775 => x"EAFFFF4C",
000776 => x"E3740001",
000777 => x"0AFFFF18",
000778 => x"E3540030",
000779 => x"0A000004",
000780 => x"E20400FF",
000781 => x"EBFFFD69",
000782 => x"E59F0490",
000783 => x"EBFFFE3A",
000784 => x"EAFFFF11",
000785 => x"E1A00004",
000786 => x"EBFFFD64",
000787 => x"EAFFFF40",
000788 => x"E1A00004",
000789 => x"EBFFFD61",
000790 => x"E59F0474",
000791 => x"EBFFFE32",
000792 => x"EBFFFD58",
000793 => x"E3700001",
000794 => x"0AFFFFFC",
000795 => x"EBFFFD55",
000796 => x"E3700001",
000797 => x"1AFFFFFC",
000798 => x"E3A05401",
000799 => x"E5950000",
000800 => x"E1A0100A",
000801 => x"E3A02008",
000802 => x"EBFFFE52",
000803 => x"E5DD0006",
000804 => x"E3500000",
000805 => x"0A000005",
000806 => x"E3A04000",
000807 => x"E2844001",
000808 => x"EBFFFD4E",
000809 => x"E7D4000A",
000810 => x"E3500000",
000811 => x"1AFFFFFA",
000812 => x"E3A00020",
000813 => x"EBFFFD49",
000814 => x"EBFFFD42",
000815 => x"E3700001",
000816 => x"1A000005",
000817 => x"E3A03401",
000818 => x"E2833E9E",
000819 => x"E2855004",
000820 => x"E2833004",
000821 => x"E1550003",
000822 => x"1AFFFFE7",
000823 => x"E59F03F4",
000824 => x"EBFFFE11",
000825 => x"EAFFFEE8",
000826 => x"E3540035",
000827 => x"0A0000AE",
000828 => x"E3540061",
000829 => x"1AFFFFCD",
000830 => x"E1A00004",
000831 => x"EBFFFD37",
000832 => x"E59F03D4",
000833 => x"EBFFFE08",
000834 => x"E59F03D0",
000835 => x"EBFFFE06",
000836 => x"E59F03CC",
000837 => x"EBFFFE04",
000838 => x"EAFFFEDB",
000839 => x"E59F03C4",
000840 => x"EBFFFE01",
000841 => x"E1A00009",
000842 => x"E3A01004",
000843 => x"E3A02000",
000844 => x"EBFFFE0B",
000845 => x"E5DD300F",
000846 => x"E3530053",
000847 => x"1A000002",
000848 => x"E5DD2010",
000849 => x"E352004D",
000850 => x"0A000004",
000851 => x"E59F0398",
000852 => x"EBFFFDF5",
000853 => x"E59F0394",
000854 => x"EBFFFDF3",
000855 => x"EAFFFECA",
000856 => x"E5DD1011",
000857 => x"E3510042",
000858 => x"1AFFFFF7",
000859 => x"E5DD0012",
000860 => x"E3500052",
000861 => x"1AFFFFF4",
000862 => x"E3A04000",
000863 => x"E5C43000",
000864 => x"E1A00000",
000865 => x"E5C42001",
000866 => x"E1A00000",
000867 => x"E5C41002",
000868 => x"E1A00000",
000869 => x"E5C40003",
000870 => x"E1A00000",
000871 => x"E241103E",
000872 => x"E1A00009",
000873 => x"E1A02004",
000874 => x"EBFFFDED",
000875 => x"E5DD300F",
000876 => x"E5C43004",
000877 => x"E5DD2010",
000878 => x"E5C42005",
000879 => x"E5DD3011",
000880 => x"E5C43006",
000881 => x"E5DD2012",
000882 => x"E1A00009",
000883 => x"E5C42007",
000884 => x"EBFFFE63",
000885 => x"E3A03CFF",
000886 => x"E28330FC",
000887 => x"E1500003",
000888 => x"E1A05000",
000889 => x"8A00009A",
000890 => x"E3700004",
000891 => x"12844008",
000892 => x"1280600B",
000893 => x"0A000006",
000894 => x"EBFFFCF2",
000895 => x"E3700001",
000896 => x"0AFFFFFC",
000897 => x"E1560004",
000898 => x"E5C40000",
000899 => x"E2844001",
000900 => x"1AFFFFF8",
000901 => x"E59F02D8",
000902 => x"EBFFFDC3",
000903 => x"E59F02D4",
000904 => x"EBFFFDC1",
000905 => x"E375000C",
000906 => x"0A00000F",
000907 => x"E3A04000",
000908 => x"E285700C",
000909 => x"E1A06004",
000910 => x"E5D45000",
000911 => x"E3A00077",
000912 => x"E1A01008",
000913 => x"E1A02006",
000914 => x"E3A03002",
000915 => x"E58D5000",
000916 => x"EBFFFD1E",
000917 => x"E3500000",
000918 => x"1AFFFFF7",
000919 => x"E2844001",
000920 => x"E1540007",
000921 => x"E1A06004",
000922 => x"1AFFFFF2",
000923 => x"E59F0288",
000924 => x"EBFFFDAD",
000925 => x"EAFFFFB6",
000926 => x"E1A00004",
000927 => x"EBFFFCD7",
000928 => x"E59F0278",
000929 => x"EBFFFDA8",
000930 => x"E59F0274",
000931 => x"EBFFFDA6",
000932 => x"E59F0270",
000933 => x"EBFFFDA4",
000934 => x"E59F026C",
000935 => x"EBFFFDA2",
000936 => x"E59F0268",
000937 => x"EBFFFDA0",
000938 => x"E59F0264",
000939 => x"EBFFFD9E",
000940 => x"E59F0260",
000941 => x"EBFFFD9C",
000942 => x"E59F025C",
000943 => x"EBFFFD9A",
000944 => x"E59F0258",
000945 => x"EBFFFD98",
000946 => x"E59F0254",
000947 => x"EBFFFD96",
000948 => x"E59F0250",
000949 => x"EBFFFD94",
000950 => x"E59F024C",
000951 => x"EBFFFD92",
000952 => x"E59F0248",
000953 => x"EBFFFD90",
000954 => x"E59F0244",
000955 => x"EBFFFD8E",
000956 => x"E59F0240",
000957 => x"EBFFFD8C",
000958 => x"E59F023C",
000959 => x"EBFFFD8A",
000960 => x"E59F0238",
000961 => x"EBFFFD88",
000962 => x"E59F0234",
000963 => x"EBFFFD86",
000964 => x"E59F0230",
000965 => x"EBFFFD84",
000966 => x"E59F022C",
000967 => x"EBFFFD82",
000968 => x"EAFFFE59",
000969 => x"E5DD3011",
000970 => x"E3530042",
000971 => x"1AFFFEE6",
000972 => x"E5DD3012",
000973 => x"E3530052",
000974 => x"1AFFFEE3",
000975 => x"E3A01004",
000976 => x"E3A02000",
000977 => x"E1A00009",
000978 => x"EBFFFD85",
000979 => x"E1A00009",
000980 => x"EBFFFE03",
000981 => x"E3A03C7F",
000982 => x"E28330F8",
000983 => x"E1500003",
000984 => x"8A00003B",
000985 => x"E2804401",
000986 => x"E2844004",
000987 => x"E3540401",
000988 => x"0A000009",
000989 => x"E3A05401",
000990 => x"E3A01004",
000991 => x"E3A02000",
000992 => x"E1A00009",
000993 => x"EBFFFD76",
000994 => x"E1A00009",
000995 => x"EBFFFDF4",
000996 => x"E4850004",
000997 => x"E1550004",
000998 => x"1AFFFFF6",
000999 => x"E59F00FC",
001000 => x"EBFFFD61",
001001 => x"EBFFFDF6",
001002 => x"EAFFFE37",
001003 => x"E1A00004",
001004 => x"EBFFFC8A",
001005 => x"E59F0194",
001006 => x"EBFFFD5B",
001007 => x"E1A00009",
001008 => x"E3A01002",
001009 => x"E3A02001",
001010 => x"EBFFFD65",
001011 => x"E1A00009",
001012 => x"E3A01002",
001013 => x"EBFFFDC7",
001014 => x"E21060FF",
001015 => x"0AFFFE89",
001016 => x"E59F016C",
001017 => x"EBFFFD50",
001018 => x"E59F0168",
001019 => x"EBFFFD4E",
001020 => x"EBFFFC74",
001021 => x"E3700001",
001022 => x"0AFFFFFC",
001023 => x"EBFFFC71",
001024 => x"E3700001",
001025 => x"1AFFFFFC",
001026 => x"E3A05000",
001027 => x"EA000001",
001028 => x"E3540000",
001029 => x"AA000011",
001030 => x"E3A0C000",
001031 => x"E1A02005",
001032 => x"E1A01006",
001033 => x"E3A03002",
001034 => x"E3A00072",
001035 => x"E58DC000",
001036 => x"EBFFFCA6",
001037 => x"E1A04000",
001038 => x"EBFFFC62",
001039 => x"E3700001",
001040 => x"E1A00004",
001041 => x"0AFFFFF1",
001042 => x"E59F010C",
001043 => x"EBFFFD36",
001044 => x"EAFFFF21",
001045 => x"E59F0104",
001046 => x"EBFFFD33",
001047 => x"EAFFFE0A",
001048 => x"EBFFFC5E",
001049 => x"E3A03801",
001050 => x"E2855001",
001051 => x"E2433001",
001052 => x"E1550003",
001053 => x"1AFFFFE7",
001054 => x"EAFFFF17",
001055 => x"0001129C",
001056 => x"000112E8",
001057 => x"00011330",
001058 => x"00011378",
001059 => x"000113C0",
001060 => x"00011408",
001061 => x"00011450",
001062 => x"000114BC",
001063 => x"000114F4",
001064 => x"00011504",
001065 => x"00011690",
001066 => x"000116F4",
001067 => x"00011DF8",
001068 => x"00011634",
001069 => x"00011670",
001070 => x"00011720",
001071 => x"00011508",
001072 => x"000115A0",
001073 => x"00011D7C",
001074 => x"00011DAC",
001075 => x"000116E0",
001076 => x"00011DD4",
001077 => x"000115C8",
001078 => x"00011610",
001079 => x"000118D0",
001080 => x"00011904",
001081 => x"00011970",
001082 => x"00011740",
001083 => x"000117E8",
001084 => x"00011DC8",
001085 => x"000117A0",
001086 => x"000117B8",
001087 => x"000117D8",
001088 => x"000119B4",
001089 => x"000119D0",
001090 => x"000119F0",
001091 => x"00011A30",
001092 => x"00011A64",
001093 => x"00011AA0",
001094 => x"00011ADC",
001095 => x"00011B00",
001096 => x"00011B3C",
001097 => x"00011B58",
001098 => x"00011B70",
001099 => x"00011BB8",
001100 => x"00011BF8",
001101 => x"00011C30",
001102 => x"00011C54",
001103 => x"00011C98",
001104 => x"00011CD8",
001105 => x"00011D04",
001106 => x"00011D30",
001107 => x"00011D54",
001108 => x"0001180C",
001109 => x"00011848",
001110 => x"00011888",
001111 => x"00011E1C",
001112 => x"0001157C",
001113 => x"E10F3000",
001114 => x"E3C330C0",
001115 => x"E129F003",
001116 => x"E1A0F00E",
001117 => x"E10F3000",
001118 => x"E38330C0",
001119 => x"E129F003",
001120 => x"E1A0F00E",
001121 => x"2030202D",
001122 => x"20626F6F",
001123 => x"74206672",
001124 => x"6F6D2063",
001125 => x"6F726520",
001126 => x"52414D20",
001127 => x"28737461",
001128 => x"72742061",
001129 => x"70706C69",
001130 => x"63617469",
001131 => x"6F6E290D",
001132 => x"0A203120",
001133 => x"2D207072",
001134 => x"6F677261",
001135 => x"6D20636F",
001136 => x"72652052",
001137 => x"414D2076",
001138 => x"69612055",
001139 => x"4152545F",
001140 => x"300D0A20",
001141 => x"32202D20",
001142 => x"636F7265",
001143 => x"2052414D",
001144 => x"2064756D",
001145 => x"700D0A00",
001146 => x"2033202D",
001147 => x"20626F6F",
001148 => x"74206672",
001149 => x"6F6D2049",
001150 => x"32432045",
001151 => x"4550524F",
001152 => x"4D0D0A20",
001153 => x"34202D20",
001154 => x"70726F67",
001155 => x"72616D20",
001156 => x"49324320",
001157 => x"45455052",
001158 => x"4F4D2076",
001159 => x"69612055",
001160 => x"4152545F",
001161 => x"300D0A20",
001162 => x"35202D20",
001163 => x"73686F77",
001164 => x"20636F6E",
001165 => x"74656E74",
001166 => x"206F6620",
001167 => x"49324320",
001168 => x"45455052",
001169 => x"4F4D0D0A",
001170 => x"00000000",
001171 => x"2061202D",
001172 => x"20617574",
001173 => x"6F6D6174",
001174 => x"69632062",
001175 => x"6F6F7420",
001176 => x"636F6E66",
001177 => x"69677572",
001178 => x"6174696F",
001179 => x"6E0D0A20",
001180 => x"68202D20",
001181 => x"68656C70",
001182 => x"0D0A2072",
001183 => x"202D2072",
001184 => x"65737461",
001185 => x"72742073",
001186 => x"79737465",
001187 => x"6D0D0A0D",
001188 => x"0A53656C",
001189 => x"6563743A",
001190 => x"20000000",
001191 => x"0D0A0D0A",
001192 => x"0D0A2B2D",
001193 => x"2D2D2D2D",
001194 => x"2D2D2D2D",
001195 => x"2D2D2D2D",
001196 => x"2D2D2D2D",
001197 => x"2D2D2D2D",
001198 => x"2D2D2D2D",
001199 => x"2D2D2D2D",
001200 => x"2D2D2D2D",
001201 => x"2D2D2D2D",
001202 => x"2D2D2D2D",
001203 => x"2D2D2D2D",
001204 => x"2D2D2D2D",
001205 => x"2D2D2D2D",
001206 => x"2D2D2D2D",
001207 => x"2D2D2D2D",
001208 => x"2D2D2D2B",
001209 => x"0D0A0000",
001210 => x"7C202020",
001211 => x"203C3C3C",
001212 => x"2053544F",
001213 => x"524D2043",
001214 => x"6F726520",
001215 => x"50726F63",
001216 => x"6573736F",
001217 => x"72205379",
001218 => x"7374656D",
001219 => x"202D2042",
001220 => x"79205374",
001221 => x"65706861",
001222 => x"6E204E6F",
001223 => x"6C74696E",
001224 => x"67203E3E",
001225 => x"3E202020",
001226 => x"207C0D0A",
001227 => x"00000000",
001228 => x"2B2D2D2D",
001229 => x"2D2D2D2D",
001230 => x"2D2D2D2D",
001231 => x"2D2D2D2D",
001232 => x"2D2D2D2D",
001233 => x"2D2D2D2D",
001234 => x"2D2D2D2D",
001235 => x"2D2D2D2D",
001236 => x"2D2D2D2D",
001237 => x"2D2D2D2D",
001238 => x"2D2D2D2D",
001239 => x"2D2D2D2D",
001240 => x"2D2D2D2D",
001241 => x"2D2D2D2D",
001242 => x"2D2D2D2D",
001243 => x"2D2D2D2D",
001244 => x"2D2B0D0A",
001245 => x"00000000",
001246 => x"7C202020",
001247 => x"20202020",
001248 => x"2020426F",
001249 => x"6F746C6F",
001250 => x"61646572",
001251 => x"20666F72",
001252 => x"2053544F",
001253 => x"524D2053",
001254 => x"6F432020",
001255 => x"20566572",
001256 => x"73696F6E",
001257 => x"3A203230",
001258 => x"31323035",
001259 => x"32342D44",
001260 => x"20202020",
001261 => x"20202020",
001262 => x"207C0D0A",
001263 => x"00000000",
001264 => x"7C202020",
001265 => x"20202020",
001266 => x"20202020",
001267 => x"20202020",
001268 => x"436F6E74",
001269 => x"6163743A",
001270 => x"2073746E",
001271 => x"6F6C7469",
001272 => x"6E674067",
001273 => x"6F6F676C",
001274 => x"656D6169",
001275 => x"6C2E636F",
001276 => x"6D202020",
001277 => x"20202020",
001278 => x"20202020",
001279 => x"20202020",
001280 => x"207C0D0A",
001281 => x"00000000",
001282 => x"2B2D2D2D",
001283 => x"2D2D2D2D",
001284 => x"2D2D2D2D",
001285 => x"2D2D2D2D",
001286 => x"2D2D2D2D",
001287 => x"2D2D2D2D",
001288 => x"2D2D2D2D",
001289 => x"2D2D2D2D",
001290 => x"2D2D2D2D",
001291 => x"2D2D2D2D",
001292 => x"2D2D2D2D",
001293 => x"2D2D2D2D",
001294 => x"2D2D2D2D",
001295 => x"2D2D2D2D",
001296 => x"2D2D2D2D",
001297 => x"2D2D2D2D",
001298 => x"2D2B0D0A",
001299 => x"0D0A0000",
001300 => x"203C2057",
001301 => x"656C636F",
001302 => x"6D652074",
001303 => x"6F207468",
001304 => x"65205354",
001305 => x"4F524D20",
001306 => x"536F4320",
001307 => x"626F6F74",
001308 => x"6C6F6164",
001309 => x"65722063",
001310 => x"6F6E736F",
001311 => x"6C652120",
001312 => x"3E0D0A20",
001313 => x"3C205365",
001314 => x"6C656374",
001315 => x"20616E20",
001316 => x"6F706572",
001317 => x"6174696F",
001318 => x"6E206672",
001319 => x"6F6D2074",
001320 => x"6865206D",
001321 => x"656E7520",
001322 => x"62656C6F",
001323 => x"77206F72",
001324 => x"20707265",
001325 => x"7373203E",
001326 => x"0D0A0000",
001327 => x"203C2074",
001328 => x"68652062",
001329 => x"6F6F7420",
001330 => x"6B657920",
001331 => x"666F7220",
001332 => x"696D6D65",
001333 => x"64696174",
001334 => x"65206170",
001335 => x"706C6963",
001336 => x"6174696F",
001337 => x"6E207374",
001338 => x"6172742E",
001339 => x"203E0D0A",
001340 => x"0D0A0000",
001341 => x"204C6F61",
001342 => x"64204164",
001343 => x"64726573",
001344 => x"733A2000",
001345 => x"0A0D0000",
001346 => x"0D0A0D0A",
001347 => x"4170706C",
001348 => x"69636174",
001349 => x"696F6E20",
001350 => x"77696C6C",
001351 => x"20737461",
001352 => x"72742061",
001353 => x"75746F6D",
001354 => x"61746963",
001355 => x"616C6C79",
001356 => x"20616674",
001357 => x"65722064",
001358 => x"6F776E6C",
001359 => x"6F61642E",
001360 => x"0D0A2D3E",
001361 => x"20576169",
001362 => x"74696E67",
001363 => x"20666F72",
001364 => x"20277374",
001365 => x"6F726D5F",
001366 => x"70726F67",
001367 => x"72616D2E",
001368 => x"62696E27",
001369 => x"20696E20",
001370 => x"62797465",
001371 => x"2D737472",
001372 => x"65616D20",
001373 => x"6D6F6465",
001374 => x"2E2E2E00",
001375 => x"20455252",
001376 => x"4F522120",
001377 => x"50726F67",
001378 => x"72616D20",
001379 => x"66696C65",
001380 => x"20746F6F",
001381 => x"20626967",
001382 => x"210D0A0D",
001383 => x"0A000000",
001384 => x"20496E76",
001385 => x"616C6964",
001386 => x"2070726F",
001387 => x"6772616D",
001388 => x"6D696E67",
001389 => x"2066696C",
001390 => x"65210D0A",
001391 => x"0D0A5365",
001392 => x"6C656374",
001393 => x"3A200000",
001394 => x"0D0A0D0A",
001395 => x"41626F72",
001396 => x"74206475",
001397 => x"6D70696E",
001398 => x"67206279",
001399 => x"20707265",
001400 => x"7373696E",
001401 => x"6720616E",
001402 => x"79206B65",
001403 => x"792E0D0A",
001404 => x"50726573",
001405 => x"7320616E",
001406 => x"79206B65",
001407 => x"7920746F",
001408 => x"20636F6E",
001409 => x"74696E75",
001410 => x"652E0D0A",
001411 => x"0D0A0000",
001412 => x"0D0A0D0A",
001413 => x"44756D70",
001414 => x"696E6720",
001415 => x"636F6D70",
001416 => x"6C657465",
001417 => x"642E0D0A",
001418 => x"0D0A5365",
001419 => x"6C656374",
001420 => x"3A200000",
001421 => x"0D0A0D0A",
001422 => x"456E7465",
001423 => x"72206465",
001424 => x"76696365",
001425 => x"20616464",
001426 => x"72657373",
001427 => x"20283278",
001428 => x"20686578",
001429 => x"5F636861",
001430 => x"72732C20",
001431 => x"73657420",
001432 => x"4C534220",
001433 => x"746F2027",
001434 => x"3027293A",
001435 => x"20000000",
001436 => x"20496E76",
001437 => x"616C6964",
001438 => x"20616464",
001439 => x"72657373",
001440 => x"210D0A0D",
001441 => x"0A53656C",
001442 => x"6563743A",
001443 => x"20000000",
001444 => x"0D0A4170",
001445 => x"706C6963",
001446 => x"6174696F",
001447 => x"6E207769",
001448 => x"6C6C2073",
001449 => x"74617274",
001450 => x"20617574",
001451 => x"6F6D6174",
001452 => x"6963616C",
001453 => x"6C792061",
001454 => x"66746572",
001455 => x"2075706C",
001456 => x"6F61642E",
001457 => x"0D0A2D3E",
001458 => x"204C6F61",
001459 => x"64696E67",
001460 => x"20626F6F",
001461 => x"7420696D",
001462 => x"6167652E",
001463 => x"2E2E0000",
001464 => x"2055706C",
001465 => x"6F616420",
001466 => x"636F6D70",
001467 => x"6C657465",
001468 => x"0D0A0000",
001469 => x"20496E76",
001470 => x"616C6964",
001471 => x"20626F6F",
001472 => x"74206465",
001473 => x"76696365",
001474 => x"206F7220",
001475 => x"66696C65",
001476 => x"210D0A0D",
001477 => x"0A53656C",
001478 => x"6563743A",
001479 => x"20000000",
001480 => x"0D0A496E",
001481 => x"76616C69",
001482 => x"64206164",
001483 => x"64726573",
001484 => x"73210D0A",
001485 => x"0D0A5365",
001486 => x"6C656374",
001487 => x"3A200000",
001488 => x"0D0A4461",
001489 => x"74612077",
001490 => x"696C6C20",
001491 => x"6F766572",
001492 => x"77726974",
001493 => x"65205241",
001494 => x"4D20636F",
001495 => x"6E74656E",
001496 => x"74210D0A",
001497 => x"2D3E2057",
001498 => x"61697469",
001499 => x"6E672066",
001500 => x"6F722027",
001501 => x"73746F72",
001502 => x"6D5F7072",
001503 => x"6F677261",
001504 => x"6D2E6269",
001505 => x"6E272069",
001506 => x"6E206279",
001507 => x"74652D73",
001508 => x"74726561",
001509 => x"6D206D6F",
001510 => x"64652E2E",
001511 => x"2E000000",
001512 => x"20446F77",
001513 => x"6E6C6F61",
001514 => x"6420636F",
001515 => x"6D706C65",
001516 => x"7465640D",
001517 => x"0A000000",
001518 => x"57726974",
001519 => x"696E6720",
001520 => x"62756666",
001521 => x"65722074",
001522 => x"6F206932",
001523 => x"63204545",
001524 => x"50524F4D",
001525 => x"2E2E2E00",
001526 => x"20436F6D",
001527 => x"706C6574",
001528 => x"65640D0A",
001529 => x"0D0A0000",
001530 => x"20496E76",
001531 => x"616C6964",
001532 => x"20626F6F",
001533 => x"74206465",
001534 => x"76696365",
001535 => x"206F7220",
001536 => x"66696C65",
001537 => x"210D0A0D",
001538 => x"0A000000",
001539 => x"0D0A0D0A",
001540 => x"456E7465",
001541 => x"72206465",
001542 => x"76696365",
001543 => x"20616464",
001544 => x"72657373",
001545 => x"20283220",
001546 => x"6865782D",
001547 => x"63686172",
001548 => x"732C2073",
001549 => x"6574204C",
001550 => x"53422074",
001551 => x"6F202730",
001552 => x"27293A20",
001553 => x"00000000",
001554 => x"0D0A0D0A",
001555 => x"41626F72",
001556 => x"74206475",
001557 => x"6D70696E",
001558 => x"67206279",
001559 => x"20707265",
001560 => x"7373696E",
001561 => x"6720616E",
001562 => x"79206B65",
001563 => x"792E2049",
001564 => x"66206E6F",
001565 => x"20646174",
001566 => x"61206973",
001567 => x"2073686F",
001568 => x"776E2C0D",
001569 => x"0A000000",
001570 => x"74686520",
001571 => x"73656C65",
001572 => x"63746564",
001573 => x"20646576",
001574 => x"69636520",
001575 => x"6973206E",
001576 => x"6F742072",
001577 => x"6573706F",
001578 => x"6E64696E",
001579 => x"672E2050",
001580 => x"72657373",
001581 => x"20616E79",
001582 => x"206B6579",
001583 => x"20746F20",
001584 => x"636F6E74",
001585 => x"696E7565",
001586 => x"2E0D0A0D",
001587 => x"0A000000",
001588 => x"0D0A0D0A",
001589 => x"4175746F",
001590 => x"6D617469",
001591 => x"6320626F",
001592 => x"6F742063",
001593 => x"6F6E6669",
001594 => x"67757261",
001595 => x"74696F6E",
001596 => x"20666F72",
001597 => x"20706F77",
001598 => x"65722D75",
001599 => x"703A0D0A",
001600 => x"00000000",
001601 => x"5B333231",
001602 => x"305D2063",
001603 => x"6F6E6669",
001604 => x"67757261",
001605 => x"74696F6E",
001606 => x"20444950",
001607 => x"20737769",
001608 => x"7463680D",
001609 => x"0A203030",
001610 => x"3030202D",
001611 => x"20537461",
001612 => x"72742062",
001613 => x"6F6F746C",
001614 => x"6F616465",
001615 => x"7220636F",
001616 => x"6E736F6C",
001617 => x"650D0A20",
001618 => x"30303031",
001619 => x"202D2041",
001620 => x"75746F6D",
001621 => x"61746963",
001622 => x"20626F6F",
001623 => x"74206672",
001624 => x"6F6D2063",
001625 => x"6F726520",
001626 => x"52414D0D",
001627 => x"0A000000",
001628 => x"20303031",
001629 => x"30202D20",
001630 => x"4175746F",
001631 => x"6D617469",
001632 => x"6320626F",
001633 => x"6F742066",
001634 => x"726F6D20",
001635 => x"49324320",
001636 => x"45455052",
001637 => x"4F4D2028",
001638 => x"41646472",
001639 => x"65737320",
001640 => x"30784130",
001641 => x"290D0A0D",
001642 => x"0A53656C",
001643 => x"6563743A",
001644 => x"20000000",
001645 => x"0D0A0D0A",
001646 => x"53544F52",
001647 => x"4D20536F",
001648 => x"4320626F",
001649 => x"6F746C6F",
001650 => x"61646572",
001651 => x"0D0A0000",
001652 => x"2730273A",
001653 => x"20457865",
001654 => x"63757465",
001655 => x"2070726F",
001656 => x"6772616D",
001657 => x"20696E20",
001658 => x"52414D2E",
001659 => x"0D0A0000",
001660 => x"2731273A",
001661 => x"20577269",
001662 => x"74652027",
001663 => x"73746F72",
001664 => x"6D5F7072",
001665 => x"6F677261",
001666 => x"6D2E6269",
001667 => x"6E272074",
001668 => x"6F207468",
001669 => x"6520636F",
001670 => x"72652773",
001671 => x"2052414D",
001672 => x"20766961",
001673 => x"20554152",
001674 => x"542E0D0A",
001675 => x"00000000",
001676 => x"2732273A",
001677 => x"20507269",
001678 => x"6E742063",
001679 => x"75727265",
001680 => x"6E742063",
001681 => x"6F6E7465",
001682 => x"6E74206F",
001683 => x"6620636F",
001684 => x"6D706C65",
001685 => x"74652063",
001686 => x"6F726520",
001687 => x"52414D2E",
001688 => x"0D0A0000",
001689 => x"2733273A",
001690 => x"204C6F61",
001691 => x"6420626F",
001692 => x"6F742069",
001693 => x"6D616765",
001694 => x"2066726F",
001695 => x"6D204545",
001696 => x"50524F4D",
001697 => x"20616E64",
001698 => x"20737461",
001699 => x"72742061",
001700 => x"70706C69",
001701 => x"63617469",
001702 => x"6F6E2E0D",
001703 => x"0A000000",
001704 => x"2734273A",
001705 => x"20577269",
001706 => x"74652027",
001707 => x"73746F72",
001708 => x"6D5F7072",
001709 => x"6F677261",
001710 => x"6D2E6269",
001711 => x"6E272074",
001712 => x"6F204932",
001713 => x"43204545",
001714 => x"50524F4D",
001715 => x"20766961",
001716 => x"20554152",
001717 => x"542E0D0A",
001718 => x"00000000",
001719 => x"2735273A",
001720 => x"20507269",
001721 => x"6E742063",
001722 => x"6F6E7465",
001723 => x"6E74206F",
001724 => x"66204932",
001725 => x"43204545",
001726 => x"50524F4D",
001727 => x"2E0D0A00",
001728 => x"2761273A",
001729 => x"2053686F",
001730 => x"77204449",
001731 => x"50207377",
001732 => x"69746368",
001733 => x"20636F6E",
001734 => x"66696775",
001735 => x"72617469",
001736 => x"6F6E7320",
001737 => x"666F7220",
001738 => x"6175746F",
001739 => x"6D617469",
001740 => x"6320626F",
001741 => x"6F742E0D",
001742 => x"0A000000",
001743 => x"2768273A",
001744 => x"2053686F",
001745 => x"77207468",
001746 => x"69732073",
001747 => x"63726565",
001748 => x"6E2E0D0A",
001749 => x"00000000",
001750 => x"2772273A",
001751 => x"20526573",
001752 => x"65742073",
001753 => x"79737465",
001754 => x"6D2E0D0A",
001755 => x"0D0A0000",
001756 => x"426F6F74",
001757 => x"20454550",
001758 => x"524F4D3A",
001759 => x"20323478",
001760 => x"786E6E6E",
001761 => x"20286C69",
001762 => x"6B652032",
001763 => x"34414136",
001764 => x"34292C20",
001765 => x"37206269",
001766 => x"74206164",
001767 => x"64726573",
001768 => x"73202B20",
001769 => x"646F6E74",
001770 => x"2D636172",
001771 => x"65206269",
001772 => x"742C0D0A",
001773 => x"00000000",
001774 => x"636F6E6E",
001775 => x"65637465",
001776 => x"6420746F",
001777 => x"20493243",
001778 => x"5F434F4E",
001779 => x"54524F4C",
001780 => x"4C45525F",
001781 => x"302C206F",
001782 => x"70657261",
001783 => x"74696E67",
001784 => x"20667265",
001785 => x"7175656E",
001786 => x"63792069",
001787 => x"73203130",
001788 => x"306B487A",
001789 => x"2C0D0A00",
001790 => x"6D617869",
001791 => x"6D756D20",
001792 => x"45455052",
001793 => x"4F4D2073",
001794 => x"697A6520",
001795 => x"3D203635",
001796 => x"35333620",
001797 => x"62797465",
001798 => x"203D3E20",
001799 => x"31362062",
001800 => x"69742061",
001801 => x"64647265",
001802 => x"73736573",
001803 => x"2C0D0A00",
001804 => x"66697865",
001805 => x"6420626F",
001806 => x"6F742064",
001807 => x"65766963",
001808 => x"65206164",
001809 => x"64726573",
001810 => x"733A2030",
001811 => x"7841300D",
001812 => x"0A0D0A00",
001813 => x"5465726D",
001814 => x"696E616C",
001815 => x"20736574",
001816 => x"75703A20",
001817 => x"39363030",
001818 => x"20626175",
001819 => x"642C2038",
001820 => x"20646174",
001821 => x"61206269",
001822 => x"74732C20",
001823 => x"6E6F2070",
001824 => x"61726974",
001825 => x"792C2031",
001826 => x"2073746F",
001827 => x"70206269",
001828 => x"740D0A0D",
001829 => x"0A000000",
001830 => x"466F7220",
001831 => x"6D6F7265",
001832 => x"20696E66",
001833 => x"6F726D61",
001834 => x"74696F6E",
001835 => x"20736565",
001836 => x"20746865",
001837 => x"2053544F",
001838 => x"524D2043",
001839 => x"6F726520",
001840 => x"2F205354",
001841 => x"4F524D20",
001842 => x"536F4320",
001843 => x"64617461",
001844 => x"73686565",
001845 => x"740D0A00",
001846 => x"68747470",
001847 => x"3A2F2F6F",
001848 => x"70656E63",
001849 => x"6F726573",
001850 => x"2E6F7267",
001851 => x"2F70726F",
001852 => x"6A656374",
001853 => x"2C73746F",
001854 => x"726D5F63",
001855 => x"6F72650D",
001856 => x"0A000000",
001857 => x"68747470",
001858 => x"3A2F2F6F",
001859 => x"70656E63",
001860 => x"6F726573",
001861 => x"2E6F7267",
001862 => x"2F70726F",
001863 => x"6A656374",
001864 => x"2C73746F",
001865 => x"726D5F73",
001866 => x"6F630D0A",
001867 => x"00000000",
001868 => x"436F6E74",
001869 => x"6163743A",
001870 => x"2073746E",
001871 => x"6F6C7469",
001872 => x"6E674067",
001873 => x"6F6F676C",
001874 => x"656D6169",
001875 => x"6C2E636F",
001876 => x"6D0D0A00",
001877 => x"28632920",
001878 => x"32303132",
001879 => x"20627920",
001880 => x"53746570",
001881 => x"68616E20",
001882 => x"4E6F6C74",
001883 => x"696E670D",
001884 => x"0A0D0A53",
001885 => x"656C6563",
001886 => x"743A2000",
001887 => x"0D0A0D0A",
001888 => x"5765276C",
001889 => x"6C207365",
001890 => x"6E642079",
001891 => x"6F752062",
001892 => x"61636B20",
001893 => x"2D20746F",
001894 => x"20746865",
001895 => x"20667574",
001896 => x"75726521",
001897 => x"2E0D0A0D",
001898 => x"0A000000",
001899 => x"202D2044",
001900 => x"6F63746F",
001901 => x"7220456D",
001902 => x"6D657420",
001903 => x"4C2E2042",
001904 => x"726F776E",
001905 => x"0D0A0D0A",
001906 => x"53656C65",
001907 => x"63743A20",
001908 => x"00000000",
001909 => x"20496E76",
001910 => x"616C6964",
001911 => x"206F7065",
001912 => x"72617469",
001913 => x"6F6E210D",
001914 => x"0A547279",
001915 => x"20616761",
001916 => x"696E3A20",
001917 => x"00000000",
001918 => x"0D0A0D0A",
001919 => x"2D3E2053",
001920 => x"74617274",
001921 => x"696E6720",
001922 => x"6170706C",
001923 => x"69636174",
001924 => x"696F6E2E",
001925 => x"2E2E0D0A",
001926 => x"0D0A0000",
001927 => x"0D0A0D0A",
001928 => x"41626F72",
001929 => x"74656421",
001930 => x"00000000",
others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;