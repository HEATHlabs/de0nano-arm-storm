-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
--				MEM_SIZE      : natural := 1024;  -- memory cells
--				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				MEM_SIZE      : natural := 2048;  -- memory cells
				LOG2_MEM_SIZE : natural := 11;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
000000 => x"EA000006",
000001 => x"EA0004AE",
000002 => x"EA0004AD",
000003 => x"EA0004AC",
000004 => x"EA0004AB",
000005 => x"EA0004AA",
000006 => x"EA0004A9",
000007 => x"EA0004A8",
000008 => x"E59F0168",
000009 => x"E10F1000",
000010 => x"E3C1107F",
000011 => x"E38110DF",
000012 => x"E129F001",
000013 => x"E1A0D000",
000014 => x"E3A00000",
000015 => x"E1A01000",
000016 => x"E1A02000",
000017 => x"E1A0B000",
000018 => x"E1A07000",
000019 => x"E59FA140",
000020 => x"E1A0E00F",
000021 => x"E1A0F00A",
000022 => x"E3A00003",
000023 => x"E13FF000",
000024 => x"E59FD098",
000025 => x"EB000209",
000026 => x"E59F1118",
000027 => x"E59F20B8",
000028 => x"E59F30B8",
000029 => x"E1520003",
000030 => x"0A000002",
000031 => x"E4924004",
000032 => x"E4814004",
000033 => x"EAFFFFFA",
000034 => x"E59F20FC",
000035 => x"E3A03000",
000036 => x"E3A04028",
000037 => x"E4823004",
000038 => x"E2544001",
000039 => x"1AFFFFFC",
000040 => x"E1A04000",
000041 => x"E38443C3",
000042 => x"E3A00000",
000043 => x"E1A0F004",
000044 => x"E92D4000",
000045 => x"E92D1FFF",
000046 => x"E3A04000",
000047 => x"E1A0500D",
000048 => x"E1A0600E",
000049 => x"E59F00CC",
000050 => x"E1A01004",
000051 => x"E4952004",
000052 => x"EB000460",
000053 => x"E354000D",
000054 => x"12844001",
000055 => x"1AFFFFF8",
000056 => x"E59F00B4",
000057 => x"E1A0100D",
000058 => x"EB00045A",
000059 => x"E59F00AC",
000060 => x"E2461004",
000061 => x"EB000457",
000062 => x"E8BD1FFF",
000063 => x"E8FD8000",
000064 => x"007FFFF8",
000065 => x"F0000020",
000066 => x"72253264",
000067 => x"20202530",
000068 => x"38780A00",
000069 => x"73702020",
000070 => x"20253038",
000071 => x"780A0070",
000072 => x"63202020",
000073 => x"25303878",
000074 => x"0A000000",
000075 => x"00010134",
000076 => x"00010184",
000077 => x"00000005",
000078 => x"54410001",
000079 => x"00000001",
000080 => x"00001000",
000081 => x"00000000",
000082 => x"00000004",
000083 => x"54410002",
000084 => x"00800000",
000085 => x"00000000",
000086 => x"00000005",
000087 => x"54410004",
000088 => x"00000001",
000089 => x"000000D0",
000090 => x"00001E00",
000091 => x"00000004",
000092 => x"54410005",
000093 => x"02700000",
000094 => x"00034000",
000095 => x"00000000",
000096 => x"00000000",
000097 => x"00000000",
000098 => x"0007C000",
000099 => x"03F01000",
000100 => x"00002100",
000101 => x"00010890",
000102 => x"00010108",
000103 => x"00010114",
000104 => x"0001011F",
000105 => x"E92D4FF0",
000106 => x"E1A04000",
000107 => x"E1A05002",
000108 => x"E1A08001",
000109 => x"E59F0170",
000110 => x"E1A01004",
000111 => x"E1A07003",
000112 => x"EB000424",
000113 => x"E59F0164",
000114 => x"E1A01005",
000115 => x"EB000421",
000116 => x"E3A03000",
000117 => x"E5853000",
000118 => x"E0846008",
000119 => x"E1A0A003",
000120 => x"E1A09008",
000121 => x"E5D61000",
000122 => x"E59F0144",
000123 => x"EB000419",
000124 => x"E5D62000",
000125 => x"E2423030",
000126 => x"E3530009",
000127 => x"E59F0134",
000128 => x"E2421041",
000129 => x"E3A0B000",
000130 => x"8A000008",
000131 => x"EB000411",
000132 => x"E5953000",
000133 => x"E1A03203",
000134 => x"E5853000",
000135 => x"E5D62000",
000136 => x"E0833002",
000137 => x"E2433030",
000138 => x"E5853000",
000139 => x"EA000022",
000140 => x"E3510005",
000141 => x"E59F0100",
000142 => x"E2423061",
000143 => x"E3A0B000",
000144 => x"8A00000A",
000145 => x"EB000403",
000146 => x"E5953000",
000147 => x"E1A03203",
000148 => x"E5853000",
000149 => x"E59F00E4",
000150 => x"EB0003FE",
000151 => x"E5D63000",
000152 => x"E5952000",
000153 => x"E0833002",
000154 => x"E2433037",
000155 => x"EA00000F",
000156 => x"E3530005",
000157 => x"E3A0B000",
000158 => x"E59F00C4",
000159 => x"8587A000",
000160 => x"83A0B001",
000161 => x"8A00000C",
000162 => x"EB0003F2",
000163 => x"E5953000",
000164 => x"E1A03203",
000165 => x"E5853000",
000166 => x"E59F00A8",
000167 => x"EB0003ED",
000168 => x"E5D63000",
000169 => x"E5952000",
000170 => x"E0833002",
000171 => x"E2433057",
000172 => x"E5853000",
000173 => x"E59F0090",
000174 => x"EB0003E6",
000175 => x"E2894001",
000176 => x"E35A0008",
000177 => x"E59F0084",
000178 => x"E2866001",
000179 => x"E1A01004",
000180 => x"E1A09004",
000181 => x"1A000005",
000182 => x"E587A000",
000183 => x"EB0003DD",
000184 => x"E5951000",
000185 => x"E59F0068",
000186 => x"EB0003DA",
000187 => x"EA000006",
000188 => x"EB0003D8",
000189 => x"E59F0058",
000190 => x"E5951000",
000191 => x"EB0003D5",
000192 => x"E35B0000",
000193 => x"E28AA001",
000194 => x"0AFFFFB5",
000195 => x"E5971000",
000196 => x"E59F0040",
000197 => x"EB0003CF",
000198 => x"E2880001",
000199 => x"E1540000",
000200 => x"D3A00000",
000201 => x"C3A00001",
000202 => x"E8BD8FF0",
000203 => x"00011E80",
000204 => x"00011E88",
000205 => x"00011E94",
000206 => x"00011EA0",
000207 => x"00011EAC",
000208 => x"00011EB8",
000209 => x"00011ED0",
000210 => x"00011EDC",
000211 => x"00011EC4",
000212 => x"00011EEC",
000213 => x"00011EF8",
000214 => x"00011F04",
000215 => x"E92D4070",
000216 => x"E24DD004",
000217 => x"E1A06002",
000218 => x"E1A0300D",
000219 => x"E1A02001",
000220 => x"E3A01002",
000221 => x"E1A04000",
000222 => x"EBFFFF89",
000223 => x"E2501000",
000224 => x"E1A0500D",
000225 => x"E1A02006",
000226 => x"E1A00004",
000227 => x"E1A0300D",
000228 => x"0A000003",
000229 => x"E59D1000",
000230 => x"E2811003",
000231 => x"EBFFFF80",
000232 => x"E1A01000",
000233 => x"E1A00001",
000234 => x"E28DD004",
000235 => x"E8BD8070",
000236 => x"E92D4010",
000237 => x"E1A04000",
000238 => x"EA000000",
000239 => x"EB0003A5",
000240 => x"E2544001",
000241 => x"E59F0004",
000242 => x"2AFFFFFB",
000243 => x"E8BD8010",
000244 => x"00011EA8",
000245 => x"E52DE004",
000246 => x"E59F00CC",
000247 => x"EB00039D",
000248 => x"E59F00C8",
000249 => x"EB00039B",
000250 => x"E3A0001D",
000251 => x"EBFFFFEF",
000252 => x"E59F00BC",
000253 => x"EB000397",
000254 => x"E59F00B8",
000255 => x"EB000395",
000256 => x"E3A00013",
000257 => x"EBFFFFE9",
000258 => x"E59F00AC",
000259 => x"EB000391",
000260 => x"E59F00A8",
000261 => x"EB00038F",
000262 => x"E59F00A4",
000263 => x"EB00038D",
000264 => x"E3A0001D",
000265 => x"EBFFFFE1",
000266 => x"E59F0098",
000267 => x"EB000389",
000268 => x"E59F0094",
000269 => x"EB000387",
000270 => x"E3A00013",
000271 => x"EBFFFFDB",
000272 => x"E59F0088",
000273 => x"EB000383",
000274 => x"E59F0084",
000275 => x"EB000381",
000276 => x"E3A00013",
000277 => x"EBFFFFD5",
000278 => x"E59F0078",
000279 => x"EB00037D",
000280 => x"E59F0074",
000281 => x"EB00037B",
000282 => x"E3A00013",
000283 => x"EBFFFFCF",
000284 => x"E59F0068",
000285 => x"EB000377",
000286 => x"E59F0064",
000287 => x"EB000375",
000288 => x"E3A0001D",
000289 => x"EBFFFFC9",
000290 => x"E59F0058",
000291 => x"EB000371",
000292 => x"E59F0054",
000293 => x"EB00036F",
000294 => x"E3A0000B",
000295 => x"EBFFFFC3",
000296 => x"E59F0048",
000297 => x"E49DE004",
000298 => x"EA00036A",
000299 => x"00011F08",
000300 => x"00011F14",
000301 => x"00011F18",
000302 => x"00011F2C",
000303 => x"00011F38",
000304 => x"00011F5C",
000305 => x"00011F88",
000306 => x"00011F8C",
000307 => x"00011FA4",
000308 => x"00011FB0",
000309 => x"00011FDC",
000310 => x"00011FE8",
000311 => x"0001200C",
000312 => x"00012018",
000313 => x"00012024",
000314 => x"00012028",
000315 => x"00012038",
000316 => x"0001204C",
000317 => x"E1A01000",
000318 => x"E5912000",
000319 => x"E59F0000",
000320 => x"EA000354",
000321 => x"0001205C",
000322 => x"E2400001",
000323 => x"E92D4010",
000324 => x"E1A04001",
000325 => x"E3500004",
000326 => x"979FF100",
000327 => x"EA000039",
000328 => x"00010534",
000329 => x"00010574",
000330 => x"00010588",
000331 => x"000105B4",
000332 => x"000105D8",
000333 => x"E59F10EC",
000334 => x"E59F00EC",
000335 => x"EB000345",
000336 => x"E3A01602",
000337 => x"E3A00505",
000338 => x"EB000153",
000339 => x"E3500602",
000340 => x"E1A04000",
000341 => x"81A01000",
000342 => x"8A000027",
000343 => x"E59F00CC",
000344 => x"EB00033C",
000345 => x"E1A01004",
000346 => x"E3A00505",
000347 => x"E8BD4010",
000348 => x"EA0001EE",
000349 => x"EBFFFF96",
000350 => x"EBFFFECC",
000351 => x"E3A00010",
000352 => x"EBFFFF8A",
000353 => x"EA000008",
000354 => x"E3A01702",
000355 => x"E59F00A0",
000356 => x"EB000330",
000357 => x"E3A00010",
000358 => x"EBFFFF84",
000359 => x"E59F0094",
000360 => x"EB00032C",
000361 => x"E3A00702",
000362 => x"EBFFFEAE",
000363 => x"E8BD4010",
000364 => x"EA000346",
000365 => x"E3A01901",
000366 => x"E59F0074",
000367 => x"EB000325",
000368 => x"E3A00010",
000369 => x"EBFFFF79",
000370 => x"E59F0068",
000371 => x"EB000321",
000372 => x"E3A00901",
000373 => x"EAFFFFF3",
000374 => x"E59F1048",
000375 => x"E59F0048",
000376 => x"EB00031C",
000377 => x"E1A00004",
000378 => x"E3A01602",
000379 => x"EB00012A",
000380 => x"E3500602",
000381 => x"98BD8010",
000382 => x"E1A01000",
000383 => x"E59F0038",
000384 => x"E8BD4010",
000385 => x"EA000313",
000386 => x"E59F0024",
000387 => x"EB000311",
000388 => x"E3A00010",
000389 => x"EBFFFF65",
000390 => x"E59F0018",
000391 => x"EB00030D",
000392 => x"E1A00004",
000393 => x"EAFFFFDF",
000394 => x"00012078",
000395 => x"00012074",
000396 => x"000120D8",
000397 => x"000120E4",
000398 => x"00011E90",
000399 => x"000120B8",
000400 => x"E92D4010",
000401 => x"E59F3238",
000402 => x"E5D0C001",
000403 => x"E1A0E000",
000404 => x"E893000F",
000405 => x"E24DD020",
000406 => x"E35C0000",
000407 => x"E1A0400D",
000408 => x"E88D000F",
000409 => x"0A000084",
000410 => x"E35C000D",
000411 => x"1A000011",
000412 => x"E5DE0000",
000413 => x"E350006C",
000414 => x"0A000005",
000415 => x"E3500073",
000416 => x"0A000006",
000417 => x"E3500068",
000418 => x"1A00000C",
000419 => x"EBFFFF50",
000420 => x"EA000079",
000421 => x"E3A00001",
000422 => x"E3A01000",
000423 => x"EA000034",
000424 => x"EBFFFE82",
000425 => x"E3A00010",
000426 => x"EBFFFF40",
000427 => x"E59F01D4",
000428 => x"EB0002E8",
000429 => x"EA000070",
000430 => x"E35C0020",
000431 => x"0A000002",
000432 => x"E59F01C4",
000433 => x"E1A0100D",
000434 => x"EA00006A",
000435 => x"E5DE3000",
000436 => x"E353006A",
000437 => x"0A00001D",
000438 => x"8A000004",
000439 => x"E3530062",
000440 => x"0A00004D",
000441 => x"E3530064",
000442 => x"1A000060",
000443 => x"EA000006",
000444 => x"E3530072",
000445 => x"0A000040",
000446 => x"E3530077",
000447 => x"0A00004F",
000448 => x"E3530070",
000449 => x"1A000059",
000450 => x"EA00001B",
000451 => x"E1A0000E",
000452 => x"E28D1010",
000453 => x"E28D2014",
000454 => x"EBFFFF0F",
000455 => x"E3500000",
000456 => x"159D4010",
000457 => x"1A000001",
000458 => x"EA000053",
000459 => x"EBFFFF70",
000460 => x"E59D3010",
000461 => x"E59D2014",
000462 => x"E0833002",
000463 => x"E1540003",
000464 => x"E1A00004",
000465 => x"E2844004",
000466 => x"3AFFFFF7",
000467 => x"EA00004A",
000468 => x"E1A0000E",
000469 => x"E3A01002",
000470 => x"E28D2010",
000471 => x"E28D3018",
000472 => x"EBFFFE8F",
000473 => x"E3500000",
000474 => x"0A000043",
000475 => x"E3A00000",
000476 => x"E59D1010",
000477 => x"EBFFFF63",
000478 => x"EA00003F",
000479 => x"E1A0000E",
000480 => x"E3A01002",
000481 => x"E28D2010",
000482 => x"E28D3018",
000483 => x"EBFFFE84",
000484 => x"E3500000",
000485 => x"0A000038",
000486 => x"E3A03000",
000487 => x"E58D3018",
000488 => x"E59D3010",
000489 => x"E4D34001",
000490 => x"E58D3010",
000491 => x"EA00000B",
000492 => x"E3540000",
000493 => x"0A000003",
000494 => x"EB0002C8",
000495 => x"E354000D",
000496 => x"E59F00C0",
000497 => x"0B0002A3",
000498 => x"E59D2010",
000499 => x"E59D3018",
000500 => x"E4D24001",
000501 => x"E2833001",
000502 => x"E58D2010",
000503 => x"E58D3018",
000504 => x"E3140080",
000505 => x"E1A00004",
000506 => x"1A000023",
000507 => x"E59D3018",
000508 => x"E3530A01",
000509 => x"3AFFFFED",
000510 => x"EA00001F",
000511 => x"E1A0000E",
000512 => x"E3A01002",
000513 => x"E28D2010",
000514 => x"E28D3018",
000515 => x"EBFFFE64",
000516 => x"E3500000",
000517 => x"0A000018",
000518 => x"EA000011",
000519 => x"E1A0000E",
000520 => x"E3A01002",
000521 => x"E28D2010",
000522 => x"E28D3018",
000523 => x"EBFFFE5C",
000524 => x"E3500000",
000525 => x"13A00005",
000526 => x"1AFFFFCC",
000527 => x"EA00000E",
000528 => x"E1A0000E",
000529 => x"E28D1010",
000530 => x"E28D201C",
000531 => x"EBFFFEC2",
000532 => x"E3500000",
000533 => x"0A000008",
000534 => x"E59D201C",
000535 => x"E59D3010",
000536 => x"E5832000",
000537 => x"E59D0010",
000538 => x"EBFFFF21",
000539 => x"EA000002",
000540 => x"E59F0014",
000541 => x"E1A0100D",
000542 => x"EB000276",
000543 => x"E28DD020",
000544 => x"E8BD8010",
000545 => x"000120F0",
000546 => x"00011E90",
000547 => x"00012074",
000548 => x"E92D41F0",
000549 => x"E3A0100C",
000550 => x"E24DD028",
000551 => x"E59F2170",
000552 => x"E59F0170",
000553 => x"EB00026B",
000554 => x"EBFFFEC9",
000555 => x"E59F0168",
000556 => x"EB000268",
000557 => x"E3A06000",
000558 => x"E1A07006",
000559 => x"E1A08006",
000560 => x"EA000001",
000561 => x"E1A06008",
000562 => x"E3A07000",
000563 => x"E3A00FFA",
000564 => x"EB00028A",
000565 => x"E2504000",
000566 => x"BAFFFFFB",
000567 => x"E354001B",
000568 => x"0A00001C",
000569 => x"E3570001",
000570 => x"0354005B",
000571 => x"13A05000",
000572 => x"03A05001",
000573 => x"03A07002",
000574 => x"0A00001D",
000575 => x"E3570002",
000576 => x"1A000038",
000577 => x"E3540041",
000578 => x"01A04005",
000579 => x"11A07005",
000580 => x"1AFFFFED",
000581 => x"EA000000",
000582 => x"EB000270",
000583 => x"E1540006",
000584 => x"E3A00008",
000585 => x"E2844001",
000586 => x"BAFFFFFA",
000587 => x"E3A04000",
000588 => x"EA000005",
000589 => x"E28D3014",
000590 => x"E7D42003",
000591 => x"E1A00002",
000592 => x"E7C4200D",
000593 => x"EB000265",
000594 => x"E2844001",
000595 => x"E1540008",
000596 => x"BAFFFFF7",
000597 => x"EAFFFFDA",
000598 => x"E3A07001",
000599 => x"EA000004",
000600 => x"E28D2028",
000601 => x"E0823006",
000602 => x"E5434028",
000603 => x"E2866001",
000604 => x"E3A07000",
000605 => x"E3560012",
000606 => x"D3A03000",
000607 => x"C3A03001",
000608 => x"E354000D",
000609 => x"03833001",
000610 => x"E3530000",
000611 => x"0AFFFFCE",
000612 => x"E3560001",
000613 => x"DA000007",
000614 => x"E3A01000",
000615 => x"E7D1200D",
000616 => x"E28D3014",
000617 => x"E7C12003",
000618 => x"E2811001",
000619 => x"E3510014",
000620 => x"1AFFFFF9",
000621 => x"E2468001",
000622 => x"E28D2028",
000623 => x"E0823006",
000624 => x"E3A04000",
000625 => x"E5434028",
000626 => x"E59F0050",
000627 => x"EB000221",
000628 => x"E1A0000D",
000629 => x"EBFFFF19",
000630 => x"E59F0044",
000631 => x"EB00021D",
000632 => x"E1A06004",
000633 => x"EAFFFFB8",
000634 => x"EB00023C",
000635 => x"E3540008",
000636 => x"13A03000",
000637 => x"03A03001",
000638 => x"E3560000",
000639 => x"D3A03000",
000640 => x"E3530000",
000641 => x"12466001",
000642 => x"11A07005",
000643 => x"1AFFFFD8",
000644 => x"EAFFFFD2",
000645 => x"00012134",
000646 => x"00012100",
000647 => x"00012140",
000648 => x"00011E90",
000649 => x"0001214C",
000650 => x"E92D4010",
000651 => x"E3A0C000",
000652 => x"E1A04000",
000653 => x"E1A0E00C",
000654 => x"E1A00001",
000655 => x"EA00000A",
000656 => x"E7DE3004",
000657 => x"E023342C",
000658 => x"E1A03083",
000659 => x"E0832001",
000660 => x"E7D31001",
000661 => x"E5D23001",
000662 => x"E1833401",
000663 => x"E023340C",
000664 => x"E1A03803",
000665 => x"E28EE001",
000666 => x"E1A0C823",
000667 => x"E15E0000",
000668 => x"E59F1008",
000669 => x"BAFFFFF1",
000670 => x"E1A0000C",
000671 => x"E8BD8010",
000672 => x"00011C80",
000673 => x"E52DE004",
000674 => x"E3A00F4B",
000675 => x"EB00021B",
000676 => x"E3500000",
000677 => x"AAFFFFFB",
000678 => x"E49DF004",
000679 => x"E92D4FF0",
000680 => x"E3A07000",
000681 => x"E24DDB01",
000682 => x"E24DD008",
000683 => x"E1A0B000",
000684 => x"E1A09001",
000685 => x"E3A0A019",
000686 => x"E3A04043",
000687 => x"E3A08001",
000688 => x"E1A06007",
000689 => x"EA000000",
000690 => x"E3A04015",
000691 => x"E3A05000",
000692 => x"E3540000",
000693 => x"11A00004",
000694 => x"1B000200",
000695 => x"E3A00FFA",
000696 => x"EB000206",
000697 => x"E3500000",
000698 => x"BA000019",
000699 => x"E3500002",
000700 => x"0A000025",
000701 => x"CA000002",
000702 => x"E3500001",
000703 => x"1A000014",
000704 => x"EA000004",
000705 => x"E3500004",
000706 => x"0A000004",
000707 => x"E3500018",
000708 => x"1A00000F",
000709 => x"EA000005",
000710 => x"E3A05080",
000711 => x"EA00001B",
000712 => x"E3A00006",
000713 => x"EB0001ED",
000714 => x"EBFFFFD5",
000715 => x"EA00007B",
000716 => x"E3A00FFA",
000717 => x"EB0001F1",
000718 => x"E3500018",
000719 => x"1A000004",
000720 => x"EBFFFFCF",
000721 => x"E3A00006",
000722 => x"EB0001E4",
000723 => x"E3E06000",
000724 => x"EA000072",
000725 => x"E2855001",
000726 => x"E3550050",
000727 => x"1AFFFFDB",
000728 => x"E3540043",
000729 => x"0AFFFFD7",
000730 => x"EBFFFFC5",
000731 => x"E3A00018",
000732 => x"EB0001DA",
000733 => x"E3A00018",
000734 => x"EB0001D8",
000735 => x"E3A00018",
000736 => x"EB0001D6",
000737 => x"E3E06001",
000738 => x"EA000064",
000739 => x"E3A05B01",
000740 => x"E3540043",
000741 => x"03A07001",
000742 => x"E1A00000",
000743 => x"E3A04000",
000744 => x"E5CD0002",
000745 => x"EA000006",
000746 => x"EB0001D4",
000747 => x"E28D3008",
000748 => x"E3500000",
000749 => x"E2433006",
000750 => x"E2844001",
000751 => x"BA000052",
000752 => x"E7C40003",
000753 => x"E3570000",
000754 => x"13A03004",
000755 => x"03A03003",
000756 => x"E0853003",
000757 => x"E1540003",
000758 => x"E3A00FFA",
000759 => x"BAFFFFF1",
000760 => x"E5DD3004",
000761 => x"E5DD2003",
000762 => x"E1E03003",
000763 => x"E20330FF",
000764 => x"E1520003",
000765 => x"1A000044",
000766 => x"E1520008",
000767 => x"0A000002",
000768 => x"E2483001",
000769 => x"E1520003",
000770 => x"1A00003F",
000771 => x"E3570000",
000772 => x"E28D4008",
000773 => x"E2444006",
000774 => x"01A01007",
000775 => x"02840003",
000776 => x"01A02001",
000777 => x"0A00000D",
000778 => x"E2840003",
000779 => x"E1A01005",
000780 => x"EBFFFF7C",
000781 => x"E0843005",
000782 => x"E5D32004",
000783 => x"E5D33003",
000784 => x"E0822403",
000785 => x"E1A02802",
000786 => x"E1500822",
000787 => x"1A00002E",
000788 => x"EA00000C",
000789 => x"E5503001",
000790 => x"E0813003",
000791 => x"E20310FF",
000792 => x"E1520005",
000793 => x"E2800001",
000794 => x"E2822001",
000795 => x"BAFFFFF8",
000796 => x"E28D2B01",
000797 => x"E2822008",
000798 => x"E0823005",
000799 => x"E5533403",
000800 => x"E1530001",
000801 => x"1A000020",
000802 => x"E5DD3003",
000803 => x"E1530008",
000804 => x"1A00000F",
000805 => x"E0663009",
000806 => x"E1550003",
000807 => x"B1A04005",
000808 => x"A1A04003",
000809 => x"E3540000",
000810 => x"DA000005",
000811 => x"E28D1008",
000812 => x"E08B0006",
000813 => x"E2411003",
000814 => x"E1A02004",
000815 => x"EB0002A0",
000816 => x"E0866004",
000817 => x"E2883001",
000818 => x"E20380FF",
000819 => x"E3A0A019",
000820 => x"EA00000B",
000821 => x"E24AA001",
000822 => x"E35A0000",
000823 => x"CA000008",
000824 => x"EBFFFF67",
000825 => x"E3A00018",
000826 => x"EB00017C",
000827 => x"E3A00018",
000828 => x"EB00017A",
000829 => x"E3A00018",
000830 => x"EB000178",
000831 => x"E3E06002",
000832 => x"EA000006",
000833 => x"E3A00006",
000834 => x"EA000001",
000835 => x"EBFFFF5C",
000836 => x"E3A00015",
000837 => x"EB000171",
000838 => x"E3A04000",
000839 => x"EAFFFF6A",
000840 => x"E1A00006",
000841 => x"E28DD008",
000842 => x"E28DDB01",
000843 => x"E8BD8FF0",
000844 => x"E92D40F0",
000845 => x"E59F1140",
000846 => x"E1A05000",
000847 => x"E3A02003",
000848 => x"E2800001",
000849 => x"EB00026A",
000850 => x"E3500000",
000851 => x"159F012C",
000852 => x"1A000006",
000853 => x"E5D52012",
000854 => x"E5D53013",
000855 => x"E1833402",
000856 => x"E3530028",
000857 => x"01A07000",
000858 => x"0A00003C",
000859 => x"E59F0110",
000860 => x"EB000138",
000861 => x"E3A00001",
000862 => x"E8BD80F0",
000863 => x"E5952020",
000864 => x"E5D5102E",
000865 => x"E5D5302F",
000866 => x"E0852002",
000867 => x"E1833401",
000868 => x"E0242397",
000869 => x"E5943004",
000870 => x"E3530001",
000871 => x"1A000018",
000872 => x"E5943014",
000873 => x"E3530000",
000874 => x"0A00002B",
000875 => x"E594300C",
000876 => x"E3530000",
000877 => x"13A06000",
000878 => x"1A00000E",
000879 => x"EA000026",
000880 => x"E5942010",
000881 => x"E0862002",
000882 => x"E0851002",
000883 => x"E5D13002",
000884 => x"E5D10003",
000885 => x"E7D5C002",
000886 => x"E1A03803",
000887 => x"E5D12001",
000888 => x"E1833C00",
000889 => x"E594E00C",
000890 => x"E183300C",
000891 => x"E1833402",
000892 => x"E78E3006",
000893 => x"E2866004",
000894 => x"E5943014",
000895 => x"E1560003",
000896 => x"3AFFFFEE",
000897 => x"E5943004",
000898 => x"E3530008",
000899 => x"1A000012",
000900 => x"E5943014",
000901 => x"E3530000",
000902 => x"0A00000F",
000903 => x"E594300C",
000904 => x"E3530000",
000905 => x"15941010",
000906 => x"1A000006",
000907 => x"EA00000A",
000908 => x"E594300C",
000909 => x"E0813003",
000910 => x"E0623003",
000911 => x"E3A02000",
000912 => x"E5832000",
000913 => x"E2811004",
000914 => x"E2842010",
000915 => x"E892000C",
000916 => x"E0823003",
000917 => x"E1510003",
000918 => x"3AFFFFF4",
000919 => x"E2877001",
000920 => x"E5D52030",
000921 => x"E5D53031",
000922 => x"E1833402",
000923 => x"E1570003",
000924 => x"3AFFFFC1",
000925 => x"E3A00000",
000926 => x"E8BD80F0",
000927 => x"00012150",
000928 => x"00012154",
000929 => x"00012170",
000930 => x"E5903000",
000931 => x"E20110FF",
000932 => x"E3530000",
000933 => x"14C31001",
000934 => x"E1A02000",
000935 => x"E1A00001",
000936 => x"15823000",
000937 => x"11A0F00E",
000938 => x"EA00010C",
000939 => x"E92D45F0",
000940 => x"E2525000",
000941 => x"E1A08000",
000942 => x"E1A07001",
000943 => x"C3A02000",
000944 => x"CA000001",
000945 => x"EA000009",
000946 => x"E2822001",
000947 => x"E7D21007",
000948 => x"E3510000",
000949 => x"1AFFFFFB",
000950 => x"E1520005",
000951 => x"A1A05001",
000952 => x"B0625005",
000953 => x"E3130002",
000954 => x"13A0A030",
000955 => x"1A000000",
000956 => x"E3A0A020",
000957 => x"E3130001",
000958 => x"13A06000",
000959 => x"01A04005",
000960 => x"0A000002",
000961 => x"EA00000A",
000962 => x"EBFFFFDE",
000963 => x"E2444001",
000964 => x"E3540000",
000965 => x"E1A00008",
000966 => x"E20A10FF",
000967 => x"CAFFFFF9",
000968 => x"E0646005",
000969 => x"E1A05004",
000970 => x"EA000001",
000971 => x"EBFFFFD5",
000972 => x"E2866001",
000973 => x"E5D73000",
000974 => x"E2531000",
000975 => x"E1A00008",
000976 => x"E2877001",
000977 => x"1AFFFFF8",
000978 => x"EA000001",
000979 => x"EBFFFFCD",
000980 => x"E2866001",
000981 => x"E3550000",
000982 => x"E1A00008",
000983 => x"E20A10FF",
000984 => x"E2455001",
000985 => x"CAFFFFF8",
000986 => x"E1A00006",
000987 => x"E8BD85F0",
000988 => x"E92D4FF0",
000989 => x"E2514000",
000990 => x"E24DD010",
000991 => x"E1A05002",
000992 => x"E1A09000",
000993 => x"E28D6034",
000994 => x"E8960C40",
000995 => x"1A000007",
000996 => x"E3A0C030",
000997 => x"E1A02006",
000998 => x"E1A0300A",
000999 => x"E1A0100D",
001000 => x"E5CDC000",
001001 => x"E5CD4001",
001002 => x"EBFFFFBF",
001003 => x"EA00003C",
001004 => x"E2533000",
001005 => x"13A03001",
001006 => x"E352000A",
001007 => x"13A03000",
001008 => x"E3530000",
001009 => x"0A000003",
001010 => x"E3540000",
001011 => x"B2644000",
001012 => x"B3A08001",
001013 => x"BA000000",
001014 => x"E3A08000",
001015 => x"E3A03000",
001016 => x"E28D700F",
001017 => x"E5CD300F",
001018 => x"EA000010",
001019 => x"E3550010",
001020 => x"0A000002",
001021 => x"EB0000CD",
001022 => x"E0030095",
001023 => x"E0633004",
001024 => x"E3530009",
001025 => x"E083200B",
001026 => x"C242303A",
001027 => x"E2833030",
001028 => x"E3550010",
001029 => x"E1A00004",
001030 => x"E1A01005",
001031 => x"E5673001",
001032 => x"01A04224",
001033 => x"0A000001",
001034 => x"EB0000C0",
001035 => x"E1A04000",
001036 => x"E3540000",
001037 => x"E1A00004",
001038 => x"E1A01005",
001039 => x"E204300F",
001040 => x"1AFFFFE9",
001041 => x"E3580000",
001042 => x"E1A02007",
001043 => x"01A04008",
001044 => x"0A00000D",
001045 => x"E3560000",
001046 => x"0A000007",
001047 => x"E31A0002",
001048 => x"0A000005",
001049 => x"E1A00009",
001050 => x"E3A0102D",
001051 => x"EBFFFF85",
001052 => x"E2466001",
001053 => x"E3A04001",
001054 => x"EA000003",
001055 => x"E3A0302D",
001056 => x"E5423001",
001057 => x"E2477001",
001058 => x"E3A04000",
001059 => x"E1A00009",
001060 => x"E1A01007",
001061 => x"E1A02006",
001062 => x"E1A0300A",
001063 => x"EBFFFF82",
001064 => x"E0840000",
001065 => x"E28DD010",
001066 => x"E8BD8FF0",
001067 => x"E92D41F0",
001068 => x"E1A07000",
001069 => x"E24DD010",
001070 => x"E1A04001",
001071 => x"E1A05002",
001072 => x"E3A06000",
001073 => x"EA00005C",
001074 => x"E3530025",
001075 => x"1A000051",
001076 => x"E5F43001",
001077 => x"E3530000",
001078 => x"0A00005A",
001079 => x"E3530025",
001080 => x"0A000050",
001081 => x"E353002D",
001082 => x"13A08000",
001083 => x"02844001",
001084 => x"03A08001",
001085 => x"EA000001",
001086 => x"E2844001",
001087 => x"E3888002",
001088 => x"E5D43000",
001089 => x"E3530030",
001090 => x"0AFFFFFA",
001091 => x"E3A0E000",
001092 => x"EA000003",
001093 => x"E3A0300A",
001094 => x"E023239E",
001095 => x"E2844001",
001096 => x"E243E030",
001097 => x"E5D42000",
001098 => x"E2423030",
001099 => x"E3530009",
001100 => x"9AFFFFF7",
001101 => x"E3520073",
001102 => x"1A000007",
001103 => x"E4953004",
001104 => x"E59F110C",
001105 => x"E3530000",
001106 => x"11A01003",
001107 => x"E1A0200E",
001108 => x"E1A03008",
001109 => x"E1A00007",
001110 => x"EA00002C",
001111 => x"E3520064",
001112 => x"1A00000A",
001113 => x"E4951004",
001114 => x"E1A00007",
001115 => x"E3A0200A",
001116 => x"E3A03001",
001117 => x"E58DE000",
001118 => x"E58D8004",
001119 => x"E3A0C061",
001120 => x"E58DC008",
001121 => x"EBFFFF79",
001122 => x"E0866000",
001123 => x"EA000029",
001124 => x"E3520078",
001125 => x"04951004",
001126 => x"01A00007",
001127 => x"03A02010",
001128 => x"0A00000E",
001129 => x"E3520058",
001130 => x"1A000007",
001131 => x"E4951004",
001132 => x"E1A00007",
001133 => x"E3A02010",
001134 => x"E3A03000",
001135 => x"E3A0C041",
001136 => x"E58DE000",
001137 => x"E58D8004",
001138 => x"EAFFFFEC",
001139 => x"E3520075",
001140 => x"1A000004",
001141 => x"E4951004",
001142 => x"E1A00007",
001143 => x"E3A0200A",
001144 => x"E3A03000",
001145 => x"EAFFFFE2",
001146 => x"E3520063",
001147 => x"1A000011",
001148 => x"E495C004",
001149 => x"E5CDC00E",
001150 => x"E3A0C000",
001151 => x"E5CDC00F",
001152 => x"E1A0200E",
001153 => x"E1A03008",
001154 => x"E1A00007",
001155 => x"E28D100E",
001156 => x"EBFFFF25",
001157 => x"EAFFFFDB",
001158 => x"E353000A",
001159 => x"01A00007",
001160 => x"03A0100D",
001161 => x"0BFFFF17",
001162 => x"E1A00007",
001163 => x"E5D41000",
001164 => x"EBFFFF14",
001165 => x"E2866001",
001166 => x"E2844001",
001167 => x"E5D43000",
001168 => x"E3530000",
001169 => x"1AFFFF9F",
001170 => x"E1A00006",
001171 => x"E28DD010",
001172 => x"E8BD81F0",
001173 => x"000121A8",
001174 => x"E92D000F",
001175 => x"E52DE004",
001176 => x"E24DD004",
001177 => x"E28D0004",
001178 => x"E3A03000",
001179 => x"E5203004",
001180 => x"E59D1008",
001181 => x"E1A0000D",
001182 => x"E28D200C",
001183 => x"EBFFFF8A",
001184 => x"E28DD004",
001185 => x"E49DE004",
001186 => x"E28DD010",
001187 => x"E1A0F00E",
001188 => x"E92D000E",
001189 => x"E52DE004",
001190 => x"E24DD004",
001191 => x"E28D3004",
001192 => x"E5230004",
001193 => x"E59D1008",
001194 => x"E1A0000D",
001195 => x"E28D200C",
001196 => x"EBFFFF7D",
001197 => x"E28DD004",
001198 => x"E49DE004",
001199 => x"E28DD00C",
001200 => x"E1A0F00E",
001201 => x"E59FB46C",
001202 => x"E58B0000",
001203 => x"EAFFFFFC",
001204 => x"E59FB460",
001205 => x"E3A0A011",
001206 => x"E58BA000",
001207 => x"EAFFFFFB",
001208 => x"E59F1454",
001209 => x"E59F3454",
001210 => x"E5932000",
001211 => x"E2022020",
001212 => x"E3520000",
001213 => x"05810000",
001214 => x"01B0F00E",
001215 => x"1AFFFFF9",
001216 => x"E59F2434",
001217 => x"E59F3434",
001218 => x"E1A01580",
001219 => x"E0811480",
001220 => x"E5930000",
001221 => x"E2100010",
001222 => x"05920000",
001223 => x"01A0F00E",
001224 => x"E2511001",
001225 => x"1AFFFFF9",
001226 => x"E3E00000",
001227 => x"E1B0F00E",
001228 => x"E92D4010",
001229 => x"E2002102",
001230 => x"E2013102",
001231 => x"E0224003",
001232 => x"E3100102",
001233 => x"11E00000",
001234 => x"12800001",
001235 => x"E3110102",
001236 => x"11E01001",
001237 => x"12811001",
001238 => x"E1A02001",
001239 => x"E1A01000",
001240 => x"E3520000",
001241 => x"0A000011",
001242 => x"E3A00000",
001243 => x"E3A03001",
001244 => x"E3530000",
001245 => x"03A03201",
001246 => x"0A000003",
001247 => x"E1520001",
001248 => x"91A02082",
001249 => x"91A03083",
001250 => x"9AFFFFF8",
001251 => x"E1510002",
001252 => x"20411002",
001253 => x"20800003",
001254 => x"E1B030A3",
001255 => x"31A020A2",
001256 => x"3AFFFFF9",
001257 => x"E3140102",
001258 => x"11E00000",
001259 => x"12800001",
001260 => x"E8FD8010",
001261 => x"E92D4070",
001262 => x"E1A06000",
001263 => x"E1862001",
001264 => x"E3120003",
001265 => x"1A00002A",
001266 => x"E8B1003C",
001267 => x"E31200FF",
001268 => x"13120CFF",
001269 => x"131208FF",
001270 => x"131204FF",
001271 => x"14862004",
001272 => x"02411004",
001273 => x"131300FF",
001274 => x"13130CFF",
001275 => x"131308FF",
001276 => x"131304FF",
001277 => x"14863004",
001278 => x"02411004",
001279 => x"131400FF",
001280 => x"13140CFF",
001281 => x"131408FF",
001282 => x"131404FF",
001283 => x"14864004",
001284 => x"02411004",
001285 => x"131500FF",
001286 => x"13150CFF",
001287 => x"131508FF",
001288 => x"131504FF",
001289 => x"14865004",
001290 => x"02411004",
001291 => x"1AFFFFE5",
001292 => x"E4913004",
001293 => x"E4C63001",
001294 => x"E21340FF",
001295 => x"08FD8070",
001296 => x"E1A03423",
001297 => x"E4C63001",
001298 => x"E21340FF",
001299 => x"08FD8070",
001300 => x"E1A03423",
001301 => x"E4C63001",
001302 => x"E21340FF",
001303 => x"08FD8070",
001304 => x"E1A03423",
001305 => x"E4C63001",
001306 => x"E21340FF",
001307 => x"08FD8070",
001308 => x"EAFFFFEE",
001309 => x"E4D13001",
001310 => x"E4C63001",
001311 => x"E3530000",
001312 => x"08FD8070",
001313 => x"E4D13001",
001314 => x"E4C63001",
001315 => x"E3530000",
001316 => x"08FD8070",
001317 => x"E4D13001",
001318 => x"E4C63001",
001319 => x"E3530000",
001320 => x"08FD8070",
001321 => x"E4D13001",
001322 => x"E4C63001",
001323 => x"E3530000",
001324 => x"08FD8070",
001325 => x"EAFFFFEE",
001326 => x"E92D41F0",
001327 => x"E1802001",
001328 => x"E3120003",
001329 => x"1A000018",
001330 => x"E8B0001C",
001331 => x"E8B100E0",
001332 => x"E1520005",
001333 => x"1A000012",
001334 => x"01530006",
001335 => x"1A00002B",
001336 => x"01540007",
001337 => x"1A000049",
001338 => x"E31200FF",
001339 => x"13120CFF",
001340 => x"131208FF",
001341 => x"131204FF",
001342 => x"131300FF",
001343 => x"13130CFF",
001344 => x"131308FF",
001345 => x"131304FF",
001346 => x"131400FF",
001347 => x"13140CFF",
001348 => x"131408FF",
001349 => x"131404FF",
001350 => x"1AFFFFEA",
001351 => x"03A00000",
001352 => x"08FD81F0",
001353 => x"E240000C",
001354 => x"E241100C",
001355 => x"E4D02001",
001356 => x"E4D13001",
001357 => x"E0324003",
001358 => x"1A00005A",
001359 => x"E4D05001",
001360 => x"E4D16001",
001361 => x"E3520000",
001362 => x"0A000054",
001363 => x"E0357006",
001364 => x"1A000054",
001365 => x"E4D02001",
001366 => x"E4D13001",
001367 => x"E3550000",
001368 => x"0A00004E",
001369 => x"E0324003",
001370 => x"1A00004E",
001371 => x"E4D05001",
001372 => x"E4D16001",
001373 => x"E3520000",
001374 => x"0A000048",
001375 => x"E0357006",
001376 => x"1A000048",
001377 => x"E3550000",
001378 => x"0A000044",
001379 => x"1AFFFFE6",
001380 => x"E31200FF",
001381 => x"13120CFF",
001382 => x"131208FF",
001383 => x"131204FF",
001384 => x"0A00003E",
001385 => x"E2400008",
001386 => x"E2411008",
001387 => x"E4D02001",
001388 => x"E4D13001",
001389 => x"E0324003",
001390 => x"1A00003A",
001391 => x"E4D05001",
001392 => x"E4D16001",
001393 => x"E3520000",
001394 => x"0A000034",
001395 => x"E0357006",
001396 => x"1A000034",
001397 => x"E4D02001",
001398 => x"E4D13001",
001399 => x"E3550000",
001400 => x"0A00002E",
001401 => x"E0324003",
001402 => x"1A00002E",
001403 => x"E4D05001",
001404 => x"E4D16001",
001405 => x"E3520000",
001406 => x"0A000028",
001407 => x"E0357006",
001408 => x"1A000028",
001409 => x"E3550000",
001410 => x"0A000024",
001411 => x"1AFFFFC6",
001412 => x"E31200FF",
001413 => x"13120CFF",
001414 => x"131208FF",
001415 => x"131204FF",
001416 => x"131300FF",
001417 => x"13130CFF",
001418 => x"131308FF",
001419 => x"131304FF",
001420 => x"0A00001A",
001421 => x"E2400004",
001422 => x"E2411004",
001423 => x"E4D02001",
001424 => x"E4D13001",
001425 => x"E0324003",
001426 => x"1A000016",
001427 => x"E4D05001",
001428 => x"E4D16001",
001429 => x"E3520000",
001430 => x"0A000010",
001431 => x"E0357006",
001432 => x"1A000010",
001433 => x"E4D02001",
001434 => x"E4D13001",
001435 => x"E3550000",
001436 => x"0A00000A",
001437 => x"E0324003",
001438 => x"1A00000A",
001439 => x"E4D05001",
001440 => x"E4D16001",
001441 => x"E3520000",
001442 => x"0A000004",
001443 => x"E0357006",
001444 => x"1A000004",
001445 => x"E3550000",
001446 => x"0A000000",
001447 => x"1AFFFFA2",
001448 => x"03A00000",
001449 => x"08FD81F0",
001450 => x"E0450006",
001451 => x"E8FD81F0",
001452 => x"E59F107C",
001453 => x"E5811000",
001454 => x"E1A0F00E",
001455 => x"E59F1070",
001456 => x"E5910000",
001457 => x"E2800801",
001458 => x"E5810000",
001459 => x"E1A0F00E",
001460 => x"E92D4010",
001461 => x"E3520000",
001462 => x"0A000004",
001463 => x"E0804002",
001464 => x"E4D13001",
001465 => x"E4C03001",
001466 => x"E1500004",
001467 => x"1AFFFFFB",
001468 => x"E8FD8010",
001469 => x"E92D4070",
001470 => x"E3520000",
001471 => x"03A00001",
001472 => x"0A00000A",
001473 => x"E3A03000",
001474 => x"E2833001",
001475 => x"E4D04001",
001476 => x"E4D15001",
001477 => x"E0546005",
001478 => x"11A00006",
001479 => x"1A000003",
001480 => x"E1530002",
001481 => x"03A00000",
001482 => x"0A000000",
001483 => x"EAFFFFF5",
001484 => x"E8FD8070",
001485 => x"07000000",
001486 => x"F0000000",
001487 => x"FFFF0200",
001488 => x"FFFF0218",
001489 => x"E3520007",
001490 => x"E92D45F0",
001491 => x"E1A0C001",
001492 => x"E1A04002",
001493 => x"E1A0A000",
001494 => x"E1A0E000",
001495 => x"83A02000",
001496 => x"8A00001E",
001497 => x"E2443001",
001498 => x"E3530006",
001499 => x"979FF103",
001500 => x"EA000140",
001501 => x"000117C8",
001502 => x"000117C0",
001503 => x"000117B8",
001504 => x"000117B0",
001505 => x"000117A8",
001506 => x"000117A0",
001507 => x"00011790",
001508 => x"E4D13001",
001509 => x"E1A0E000",
001510 => x"E4CE3001",
001511 => x"E1A0C001",
001512 => x"E4DC3001",
001513 => x"E4CE3001",
001514 => x"E4DC3001",
001515 => x"E4CE3001",
001516 => x"E4DC3001",
001517 => x"E4CE3001",
001518 => x"E4DC3001",
001519 => x"E4CE3001",
001520 => x"E4DC3001",
001521 => x"E4CE3001",
001522 => x"E5DC3000",
001523 => x"E5CE3000",
001524 => x"EA000128",
001525 => x"E7D23001",
001526 => x"E7C2300A",
001527 => x"E2822001",
001528 => x"E08AE002",
001529 => x"E31E0003",
001530 => x"1AFFFFF9",
001531 => x"E0811002",
001532 => x"E2013003",
001533 => x"E0626004",
001534 => x"E3530003",
001535 => x"979FF103",
001536 => x"EA00011B",
001537 => x"00011814",
001538 => x"000118E4",
001539 => x"000119F4",
001540 => x"00011B04",
001541 => x"E1A02126",
001542 => x"E3A0C000",
001543 => x"EA000003",
001544 => x"E79C3001",
001545 => x"E2422001",
001546 => x"E78C300E",
001547 => x"E28CC004",
001548 => x"E3120007",
001549 => x"1AFFFFF9",
001550 => x"E08E500C",
001551 => x"E081100C",
001552 => x"E1A021A2",
001553 => x"E1A0E005",
001554 => x"E1A0C001",
001555 => x"E1A04002",
001556 => x"EA00000F",
001557 => x"E51C3020",
001558 => x"E50E3020",
001559 => x"E51C301C",
001560 => x"E50E301C",
001561 => x"E51C3018",
001562 => x"E50E3018",
001563 => x"E51C3014",
001564 => x"E50E3014",
001565 => x"E51C3010",
001566 => x"E50E3010",
001567 => x"E51C300C",
001568 => x"E50E300C",
001569 => x"E51C3008",
001570 => x"E50E3008",
001571 => x"E51C3004",
001572 => x"E50E3004",
001573 => x"E2444001",
001574 => x"E3740001",
001575 => x"E28EE020",
001576 => x"E28CC020",
001577 => x"1AFFFFEA",
001578 => x"E2063003",
001579 => x"E1A02282",
001580 => x"E2433001",
001581 => x"E085C002",
001582 => x"E0811002",
001583 => x"E3530006",
001584 => x"979FF103",
001585 => x"EA0000EB",
001586 => x"00011C68",
001587 => x"00011C60",
001588 => x"00011C58",
001589 => x"00011C50",
001590 => x"00011C48",
001591 => x"00011C40",
001592 => x"00011C38",
001593 => x"E3C10003",
001594 => x"E5904000",
001595 => x"E3CE1003",
001596 => x"E1A0C126",
001597 => x"E1A02001",
001598 => x"EA000003",
001599 => x"E7954003",
001600 => x"E18E3C04",
001601 => x"E5023004",
001602 => x"E24CC001",
001603 => x"E2822004",
001604 => x"E31C0007",
001605 => x"E2615000",
001606 => x"E1A0E424",
001607 => x"E0803002",
001608 => x"1AFFFFF5",
001609 => x"E0613000",
001610 => x"E0837002",
001611 => x"E1A001AC",
001612 => x"E2428004",
001613 => x"E1A0E008",
001614 => x"E1A0C007",
001615 => x"E1A05000",
001616 => x"EA00001F",
001617 => x"E51C2020",
001618 => x"E1A03C02",
001619 => x"E1833424",
001620 => x"E50E3020",
001621 => x"E51C101C",
001622 => x"E1A03C01",
001623 => x"E1833422",
001624 => x"E50E301C",
001625 => x"E51C2018",
001626 => x"E1A03C02",
001627 => x"E1833421",
001628 => x"E50E3018",
001629 => x"E51C1014",
001630 => x"E1A03C01",
001631 => x"E1833422",
001632 => x"E50E3014",
001633 => x"E51C2010",
001634 => x"E1A03C02",
001635 => x"E1833421",
001636 => x"E50E3010",
001637 => x"E51C100C",
001638 => x"E1A03C01",
001639 => x"E1833422",
001640 => x"E50E300C",
001641 => x"E51C2008",
001642 => x"E1A03C02",
001643 => x"E1833421",
001644 => x"E50E3008",
001645 => x"E51C4004",
001646 => x"E1A03C04",
001647 => x"E1833422",
001648 => x"E50E3004",
001649 => x"E2455001",
001650 => x"E3750001",
001651 => x"E28EE020",
001652 => x"E28CC020",
001653 => x"1AFFFFDA",
001654 => x"E1A03280",
001655 => x"E2062003",
001656 => x"E0871003",
001657 => x"E2422001",
001658 => x"E088C003",
001659 => x"E2411003",
001660 => x"EA000086",
001661 => x"E3C10003",
001662 => x"E5904000",
001663 => x"E3CE1003",
001664 => x"E1A0C126",
001665 => x"E1A02001",
001666 => x"EA000003",
001667 => x"E7954003",
001668 => x"E18E3804",
001669 => x"E5023004",
001670 => x"E24CC001",
001671 => x"E2822004",
001672 => x"E31C0007",
001673 => x"E2615000",
001674 => x"E1A0E824",
001675 => x"E0803002",
001676 => x"1AFFFFF5",
001677 => x"E0613000",
001678 => x"E0837002",
001679 => x"E1A001AC",
001680 => x"E2428004",
001681 => x"E1A0E008",
001682 => x"E1A0C007",
001683 => x"E1A05000",
001684 => x"EA00001F",
001685 => x"E51C2020",
001686 => x"E1A03802",
001687 => x"E1833824",
001688 => x"E50E3020",
001689 => x"E51C101C",
001690 => x"E1A03801",
001691 => x"E1833822",
001692 => x"E50E301C",
001693 => x"E51C2018",
001694 => x"E1A03802",
001695 => x"E1833821",
001696 => x"E50E3018",
001697 => x"E51C1014",
001698 => x"E1A03801",
001699 => x"E1833822",
001700 => x"E50E3014",
001701 => x"E51C2010",
001702 => x"E1A03802",
001703 => x"E1833821",
001704 => x"E50E3010",
001705 => x"E51C100C",
001706 => x"E1A03801",
001707 => x"E1833822",
001708 => x"E50E300C",
001709 => x"E51C2008",
001710 => x"E1A03802",
001711 => x"E1833821",
001712 => x"E50E3008",
001713 => x"E51C4004",
001714 => x"E1A03804",
001715 => x"E1833822",
001716 => x"E50E3004",
001717 => x"E2455001",
001718 => x"E3750001",
001719 => x"E28EE020",
001720 => x"E28CC020",
001721 => x"1AFFFFDA",
001722 => x"E1A03280",
001723 => x"E2062003",
001724 => x"E0871003",
001725 => x"E2422001",
001726 => x"E088C003",
001727 => x"E2411002",
001728 => x"EA000042",
001729 => x"E3C10003",
001730 => x"E5904000",
001731 => x"E3CE1003",
001732 => x"E1A0C126",
001733 => x"E1A02001",
001734 => x"EA000003",
001735 => x"E7954003",
001736 => x"E18E3404",
001737 => x"E5023004",
001738 => x"E24CC001",
001739 => x"E2822004",
001740 => x"E31C0007",
001741 => x"E2615000",
001742 => x"E1A0EC24",
001743 => x"E0803002",
001744 => x"1AFFFFF5",
001745 => x"E0613000",
001746 => x"E0837002",
001747 => x"E1A001AC",
001748 => x"E2428004",
001749 => x"E1A0E008",
001750 => x"E1A0C007",
001751 => x"E1A05000",
001752 => x"EA00001F",
001753 => x"E51C2020",
001754 => x"E1A03402",
001755 => x"E1833C24",
001756 => x"E50E3020",
001757 => x"E51C101C",
001758 => x"E1A03401",
001759 => x"E1833C22",
001760 => x"E50E301C",
001761 => x"E51C2018",
001762 => x"E1A03402",
001763 => x"E1833C21",
001764 => x"E50E3018",
001765 => x"E51C1014",
001766 => x"E1A03401",
001767 => x"E1833C22",
001768 => x"E50E3014",
001769 => x"E51C2010",
001770 => x"E1A03402",
001771 => x"E1833C21",
001772 => x"E50E3010",
001773 => x"E51C100C",
001774 => x"E1A03401",
001775 => x"E1833C22",
001776 => x"E50E300C",
001777 => x"E51C2008",
001778 => x"E1A03402",
001779 => x"E1833C21",
001780 => x"E50E3008",
001781 => x"E51C4004",
001782 => x"E1A03404",
001783 => x"E1833C22",
001784 => x"E50E3004",
001785 => x"E2455001",
001786 => x"E3750001",
001787 => x"E28EE020",
001788 => x"E28CC020",
001789 => x"1AFFFFDA",
001790 => x"E1A03280",
001791 => x"E2062003",
001792 => x"E0871003",
001793 => x"E2422001",
001794 => x"E088C003",
001795 => x"E2411001",
001796 => x"E3520006",
001797 => x"979FF102",
001798 => x"EA000016",
001799 => x"00011C68",
001800 => x"00011C60",
001801 => x"00011C58",
001802 => x"00011C50",
001803 => x"00011C48",
001804 => x"00011C40",
001805 => x"00011C38",
001806 => x"E4D13001",
001807 => x"E4CC3001",
001808 => x"E4D13001",
001809 => x"E4CC3001",
001810 => x"E4D13001",
001811 => x"E4CC3001",
001812 => x"E4D13001",
001813 => x"E4CC3001",
001814 => x"E4D13001",
001815 => x"E4CC3001",
001816 => x"E4D13001",
001817 => x"E4CC3001",
001818 => x"E5D13000",
001819 => x"E5CC3000",
001820 => x"EA000000",
001821 => x"E8BD85F0",
001822 => x"E1A0000A",
001823 => x"E8BD85F0",
001824 => x"00001021",
001825 => x"20423063",
001826 => x"408450A5",
001827 => x"60C670E7",
001828 => x"81089129",
001829 => x"A14AB16B",
001830 => x"C18CD1AD",
001831 => x"E1CEF1EF",
001832 => x"12310210",
001833 => x"32732252",
001834 => x"52B54294",
001835 => x"72F762D6",
001836 => x"93398318",
001837 => x"B37BA35A",
001838 => x"D3BDC39C",
001839 => x"F3FFE3DE",
001840 => x"24623443",
001841 => x"04201401",
001842 => x"64E674C7",
001843 => x"44A45485",
001844 => x"A56AB54B",
001845 => x"85289509",
001846 => x"E5EEF5CF",
001847 => x"C5ACD58D",
001848 => x"36532672",
001849 => x"16110630",
001850 => x"76D766F6",
001851 => x"569546B4",
001852 => x"B75BA77A",
001853 => x"97198738",
001854 => x"F7DFE7FE",
001855 => x"D79DC7BC",
001856 => x"48C458E5",
001857 => x"688678A7",
001858 => x"08401861",
001859 => x"28023823",
001860 => x"C9CCD9ED",
001861 => x"E98EF9AF",
001862 => x"89489969",
001863 => x"A90AB92B",
001864 => x"5AF54AD4",
001865 => x"7AB76A96",
001866 => x"1A710A50",
001867 => x"3A332A12",
001868 => x"DBFDCBDC",
001869 => x"FBBFEB9E",
001870 => x"9B798B58",
001871 => x"BB3BAB1A",
001872 => x"6CA67C87",
001873 => x"4CE45CC5",
001874 => x"2C223C03",
001875 => x"0C601C41",
001876 => x"EDAEFD8F",
001877 => x"CDECDDCD",
001878 => x"AD2ABD0B",
001879 => x"8D689D49",
001880 => x"7E976EB6",
001881 => x"5ED54EF4",
001882 => x"3E132E32",
001883 => x"1E510E70",
001884 => x"FF9FEFBE",
001885 => x"DFDDCFFC",
001886 => x"BF1BAF3A",
001887 => x"9F598F78",
001888 => x"918881A9",
001889 => x"B1CAA1EB",
001890 => x"D10CC12D",
001891 => x"F14EE16F",
001892 => x"108000A1",
001893 => x"30C220E3",
001894 => x"50044025",
001895 => x"70466067",
001896 => x"83B99398",
001897 => x"A3FBB3DA",
001898 => x"C33DD31C",
001899 => x"E37FF35E",
001900 => x"02B11290",
001901 => x"22F332D2",
001902 => x"42355214",
001903 => x"62777256",
001904 => x"B5EAA5CB",
001905 => x"95A88589",
001906 => x"F56EE54F",
001907 => x"D52CC50D",
001908 => x"34E224C3",
001909 => x"14A00481",
001910 => x"74666447",
001911 => x"54244405",
001912 => x"A7DBB7FA",
001913 => x"879997B8",
001914 => x"E75FF77E",
001915 => x"C71DD73C",
001916 => x"26D336F2",
001917 => x"069116B0",
001918 => x"66577676",
001919 => x"46155634",
001920 => x"D94CC96D",
001921 => x"F90EE92F",
001922 => x"99C889E9",
001923 => x"B98AA9AB",
001924 => x"58444865",
001925 => x"78066827",
001926 => x"18C008E1",
001927 => x"388228A3",
001928 => x"CB7DDB5C",
001929 => x"EB3FFB1E",
001930 => x"8BF99BD8",
001931 => x"ABBBBB9A",
001932 => x"4A755A54",
001933 => x"6A377A16",
001934 => x"0AF11AD0",
001935 => x"2AB33A92",
001936 => x"FD2EED0F",
001937 => x"DD6CCD4D",
001938 => x"BDAAAD8B",
001939 => x"9DE88DC9",
001940 => x"7C266C07",
001941 => x"5C644C45",
001942 => x"3CA22C83",
001943 => x"1CE00CC1",
001944 => x"EF1FFF3E",
001945 => x"CF5DDF7C",
001946 => x"AF9BBFBA",
001947 => x"8FD99FF8",
001948 => x"6E177E36",
001949 => x"4E555E74",
001950 => x"2E933EB2",
001951 => x"0ED11EF0",
001952 => x"2573200A",
001953 => x"00000000",
001954 => x"61646472",
001955 => x"20257820",
001956 => x"0A000000",
001957 => x"63686172",
001958 => x"3A202563",
001959 => x"20000000",
001960 => x"30207468",
001961 => x"72752039",
001962 => x"20000000",
001963 => x"41207468",
001964 => x"72752046",
001965 => x"20000000",
001966 => x"73686966",
001967 => x"74206164",
001968 => x"64722000",
001969 => x"696E6372",
001970 => x"20616464",
001971 => x"72200000",
001972 => x"61207468",
001973 => x"72752066",
001974 => x"20000000",
001975 => x"73686966",
001976 => x"74206164",
001977 => x"64726573",
001978 => x"73200000",
001979 => x"63706F73",
001980 => x"3A257820",
001981 => x"00000000",
001982 => x"61646472",
001983 => x"3A25780A",
001984 => x"00000000",
001985 => x"25692000",
001986 => x"436F6D6D",
001987 => x"616E6473",
001988 => x"0A000000",
001989 => x"6C000000",
001990 => x"3A204C6F",
001991 => x"61642065",
001992 => x"6C662066",
001993 => x"696C650A",
001994 => x"00000000",
001995 => x"62203C61",
001996 => x"64647265",
001997 => x"73733E00",
001998 => x"3A204C6F",
001999 => x"61642062",
002000 => x"696E6172",
002001 => x"79206669",
002002 => x"6C652074",
002003 => x"6F203C61",
002004 => x"64647265",
002005 => x"73733E0A",
002006 => x"00000000",
002007 => x"64203C73",
002008 => x"74617274",
002009 => x"20616464",
002010 => x"72657373",
002011 => x"3E203C6E",
002012 => x"756D2062",
002013 => x"79746573",
002014 => x"3E203A20",
002015 => x"44756D70",
002016 => x"206D656D",
002017 => x"0A000000",
002018 => x"68000000",
002019 => x"3A205072",
002020 => x"696E7420",
002021 => x"68656C70",
002022 => x"206D6573",
002023 => x"73616765",
002024 => x"0A000000",
002025 => x"6A203C61",
002026 => x"64647265",
002027 => x"73733E00",
002028 => x"3A204578",
002029 => x"65637574",
002030 => x"65206C6F",
002031 => x"61646564",
002032 => x"20656C66",
002033 => x"2C206A75",
002034 => x"6D70696E",
002035 => x"6720746F",
002036 => x"203C6164",
002037 => x"64726573",
002038 => x"733E0A00",
002039 => x"70203C61",
002040 => x"64647265",
002041 => x"73733E00",
002042 => x"3A205072",
002043 => x"696E7420",
002044 => x"61736369",
002045 => x"69206D65",
002046 => x"6D20756E",
002047 => x"74696C20",
002048 => x"66697273",
002049 => x"7420300A",
002050 => x"00000000",
002051 => x"72203C61",
002052 => x"64647265",
002053 => x"73733E00",
002054 => x"3A205265",
002055 => x"6164206D",
002056 => x"656D0A00",
002057 => x"73000000",
002058 => x"3A20436F",
002059 => x"72652073",
002060 => x"74617475",
002061 => x"730A0000",
002062 => x"77203C61",
002063 => x"64647265",
002064 => x"73733E20",
002065 => x"3C76616C",
002066 => x"75653E00",
002067 => x"3A205772",
002068 => x"69746520",
002069 => x"6D656D0A",
002070 => x"00000000",
002071 => x"6D656D20",
002072 => x"30782530",
002073 => x"3878203D",
002074 => x"20307825",
002075 => x"3038780A",
002076 => x"00000000",
002077 => x"25730A00",
002078 => x"53656E64",
002079 => x"2066696C",
002080 => x"6520772F",
002081 => x"20314B20",
002082 => x"586D6F64",
002083 => x"656D2070",
002084 => x"726F746F",
002085 => x"636F6C20",
002086 => x"66726F6D",
002087 => x"20746572",
002088 => x"6D696E61",
002089 => x"6C20656D",
002090 => x"756C6174",
002091 => x"6F72206E",
002092 => x"6F772E2E",
002093 => x"2E000000",
002094 => x"586D6F64",
002095 => x"656D2065",
002096 => x"72726F72",
002097 => x"2066696C",
002098 => x"65207369",
002099 => x"7A652030",
002100 => x"78257820",
002101 => x"0A000000",
002102 => x"0A656C66",
002103 => x"2073706C",
002104 => x"69740A00",
002105 => x"6A203078",
002106 => x"25303878",
002107 => x"0A000000",
002108 => x"496E7661",
002109 => x"6C696420",
002110 => x"636F6D6D",
002111 => x"616E6400",
002112 => x"2563416D",
002113 => x"62657220",
002114 => x"426F6F74",
002115 => x"204C6F61",
002116 => x"64657220",
002117 => x"77697468",
002118 => x"20444530",
002119 => x"2D4E414E",
002120 => x"4F203332",
002121 => x"4D422073",
002122 => x"7570706F",
002123 => x"72747625",
002124 => x"730A0000",
002125 => x"32303135",
002126 => x"2D31302D",
002127 => x"30330000",
002128 => x"52656164",
002129 => x"790A3E20",
002130 => x"00000000",
002131 => x"3E200000",
002132 => x"454C4600",
002133 => x"4552524F",
002134 => x"523A204E",
002135 => x"6F742061",
002136 => x"6E20454C",
002137 => x"46206669",
002138 => x"6C652E0A",
002139 => x"00000000",
002140 => x"4552524F",
002141 => x"523A2045",
002142 => x"4C462066",
002143 => x"696C6520",
002144 => x"6E6F7420",
002145 => x"74617267",
002146 => x"65747469",
002147 => x"6E672063",
002148 => x"6F727265",
002149 => x"63742070",
002150 => x"726F6365",
002151 => x"73736F72",
002152 => x"20747970",
002153 => x"650A0000",
002154 => x"286E756C",
002155 => x"6C290000",
others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;