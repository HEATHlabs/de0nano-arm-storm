-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
--				MEM_SIZE      : natural := 1024;  -- memory cells
--				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				MEM_SIZE      : natural := 2048;  -- memory cells
				LOG2_MEM_SIZE : natural := 11;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
000000 => x"EA000006",
000001 => x"EA00049F",
000002 => x"EA00049E",
000003 => x"EA00049D",
000004 => x"EA00049C",
000005 => x"EA00049B",
000006 => x"EA00049A",
000007 => x"EA000499",
000008 => x"E59F0168",
000009 => x"E10F1000",
000010 => x"E3C1107F",
000011 => x"E38110DF",
000012 => x"E129F001",
000013 => x"E1A0D000",
000014 => x"E3A00000",
000015 => x"E1A01000",
000016 => x"E1A02000",
000017 => x"E1A0B000",
000018 => x"E1A07000",
000019 => x"E59FA140",
000020 => x"E1A0E00F",
000021 => x"E1A0F00A",
000022 => x"E3A00003",
000023 => x"E13FF000",
000024 => x"E59FD098",
000025 => x"EB0001FA",
000026 => x"E59F1118",
000027 => x"E59F20B8",
000028 => x"E59F30B8",
000029 => x"E1520003",
000030 => x"0A000002",
000031 => x"E4924004",
000032 => x"E4814004",
000033 => x"EAFFFFFA",
000034 => x"E59F20FC",
000035 => x"E3A03000",
000036 => x"E3A04028",
000037 => x"E4823004",
000038 => x"E2544001",
000039 => x"1AFFFFFC",
000040 => x"E1A04000",
000041 => x"E38443C3",
000042 => x"E3A00000",
000043 => x"E1A0F004",
000044 => x"E92D4000",
000045 => x"E92D1FFF",
000046 => x"E3A04000",
000047 => x"E1A0500D",
000048 => x"E1A0600E",
000049 => x"E59F00CC",
000050 => x"E1A01004",
000051 => x"E4952004",
000052 => x"EB000451",
000053 => x"E354000D",
000054 => x"12844001",
000055 => x"1AFFFFF8",
000056 => x"E59F00B4",
000057 => x"E1A0100D",
000058 => x"EB00044B",
000059 => x"E59F00AC",
000060 => x"E2461004",
000061 => x"EB000448",
000062 => x"E8BD1FFF",
000063 => x"E8FD8000",
000064 => x"007FFFF8",
000065 => x"F0000020",
000066 => x"72253264",
000067 => x"20202530",
000068 => x"38780A00",
000069 => x"73702020",
000070 => x"20253038",
000071 => x"780A0070",
000072 => x"63202020",
000073 => x"25303878",
000074 => x"0A000000",
000075 => x"00010134",
000076 => x"00010184",
000077 => x"00000005",
000078 => x"54410001",
000079 => x"00000001",
000080 => x"00001000",
000081 => x"00000000",
000082 => x"00000004",
000083 => x"54410002",
000084 => x"00800000",
000085 => x"00000000",
000086 => x"00000005",
000087 => x"54410004",
000088 => x"00000001",
000089 => x"000000D0",
000090 => x"00001E00",
000091 => x"00000004",
000092 => x"54410005",
000093 => x"02700000",
000094 => x"00034000",
000095 => x"00000000",
000096 => x"00000000",
000097 => x"00000000",
000098 => x"0007C000",
000099 => x"03F01000",
000100 => x"00002100",
000101 => x"00010854",
000102 => x"00010108",
000103 => x"00010114",
000104 => x"0001011F",
000105 => x"E92D4FF0",
000106 => x"E1A04000",
000107 => x"E1A08001",
000108 => x"E59F0148",
000109 => x"E1A01004",
000110 => x"E1A05002",
000111 => x"E1A07003",
000112 => x"EB000415",
000113 => x"E3A03000",
000114 => x"E5853000",
000115 => x"E0846008",
000116 => x"E1A0A003",
000117 => x"E1A09008",
000118 => x"E5D61000",
000119 => x"E59F0120",
000120 => x"EB00040D",
000121 => x"E5D62000",
000122 => x"E2423030",
000123 => x"E3530009",
000124 => x"E59F0110",
000125 => x"E2421041",
000126 => x"E3A0B000",
000127 => x"8A000007",
000128 => x"EB000405",
000129 => x"E5953000",
000130 => x"E1A03203",
000131 => x"E5853000",
000132 => x"E5D62000",
000133 => x"E0833002",
000134 => x"E2433030",
000135 => x"EA00000B",
000136 => x"E3510005",
000137 => x"E59F00E0",
000138 => x"E2423061",
000139 => x"E3A0B000",
000140 => x"8A000008",
000141 => x"EB0003F8",
000142 => x"E5953000",
000143 => x"E1A03203",
000144 => x"E5853000",
000145 => x"E5D62000",
000146 => x"E0833002",
000147 => x"E2433037",
000148 => x"E5853000",
000149 => x"EA00000D",
000150 => x"E3530005",
000151 => x"E3A0B000",
000152 => x"E59F00A8",
000153 => x"8587A000",
000154 => x"83A0B001",
000155 => x"8A000007",
000156 => x"EB0003E9",
000157 => x"E5953000",
000158 => x"E1A03203",
000159 => x"E5853000",
000160 => x"E5D62000",
000161 => x"E0833002",
000162 => x"E2433057",
000163 => x"EAFFFFEF",
000164 => x"E2894001",
000165 => x"E35A0008",
000166 => x"E59F0074",
000167 => x"E2866001",
000168 => x"E1A01004",
000169 => x"E1A09004",
000170 => x"1A000005",
000171 => x"E587A000",
000172 => x"EB0003D9",
000173 => x"E5951000",
000174 => x"E59F0058",
000175 => x"EB0003D6",
000176 => x"EA000006",
000177 => x"EB0003D4",
000178 => x"E59F0048",
000179 => x"E5951000",
000180 => x"EB0003D1",
000181 => x"E35B0000",
000182 => x"E28AA001",
000183 => x"0AFFFFBD",
000184 => x"E5971000",
000185 => x"E59F0030",
000186 => x"EB0003CB",
000187 => x"E2880001",
000188 => x"E1540000",
000189 => x"D3A00000",
000190 => x"C3A00001",
000191 => x"E8BD8FF0",
000192 => x"00011E44",
000193 => x"00011E4C",
000194 => x"00011E58",
000195 => x"00011E64",
000196 => x"00011E70",
000197 => x"00011E7C",
000198 => x"00011E88",
000199 => x"00011E94",
000200 => x"E92D4070",
000201 => x"E24DD004",
000202 => x"E1A06002",
000203 => x"E1A0300D",
000204 => x"E1A02001",
000205 => x"E3A01002",
000206 => x"E1A04000",
000207 => x"EBFFFF98",
000208 => x"E2501000",
000209 => x"E1A0500D",
000210 => x"E1A02006",
000211 => x"E1A00004",
000212 => x"E1A0300D",
000213 => x"0A000003",
000214 => x"E59D1000",
000215 => x"E2811003",
000216 => x"EBFFFF8F",
000217 => x"E1A01000",
000218 => x"E1A00001",
000219 => x"E28DD004",
000220 => x"E8BD8070",
000221 => x"E92D4010",
000222 => x"E1A04000",
000223 => x"EA000000",
000224 => x"EB0003A5",
000225 => x"E2544001",
000226 => x"E59F0004",
000227 => x"2AFFFFFB",
000228 => x"E8BD8010",
000229 => x"00011E54",
000230 => x"E52DE004",
000231 => x"E59F00CC",
000232 => x"EB00039D",
000233 => x"E59F00C8",
000234 => x"EB00039B",
000235 => x"E3A0001D",
000236 => x"EBFFFFEF",
000237 => x"E59F00BC",
000238 => x"EB000397",
000239 => x"E59F00B8",
000240 => x"EB000395",
000241 => x"E3A00013",
000242 => x"EBFFFFE9",
000243 => x"E59F00AC",
000244 => x"EB000391",
000245 => x"E59F00A8",
000246 => x"EB00038F",
000247 => x"E59F00A4",
000248 => x"EB00038D",
000249 => x"E3A0001D",
000250 => x"EBFFFFE1",
000251 => x"E59F0098",
000252 => x"EB000389",
000253 => x"E59F0094",
000254 => x"EB000387",
000255 => x"E3A00013",
000256 => x"EBFFFFDB",
000257 => x"E59F0088",
000258 => x"EB000383",
000259 => x"E59F0084",
000260 => x"EB000381",
000261 => x"E3A00013",
000262 => x"EBFFFFD5",
000263 => x"E59F0078",
000264 => x"EB00037D",
000265 => x"E59F0074",
000266 => x"EB00037B",
000267 => x"E3A00013",
000268 => x"EBFFFFCF",
000269 => x"E59F0068",
000270 => x"EB000377",
000271 => x"E59F0064",
000272 => x"EB000375",
000273 => x"E3A0001D",
000274 => x"EBFFFFC9",
000275 => x"E59F0058",
000276 => x"EB000371",
000277 => x"E59F0054",
000278 => x"EB00036F",
000279 => x"E3A0000B",
000280 => x"EBFFFFC3",
000281 => x"E59F0048",
000282 => x"E49DE004",
000283 => x"EA00036A",
000284 => x"00011E98",
000285 => x"00011EA4",
000286 => x"00011EA8",
000287 => x"00011EBC",
000288 => x"00011EC8",
000289 => x"00011EEC",
000290 => x"00011F18",
000291 => x"00011F1C",
000292 => x"00011F34",
000293 => x"00011F40",
000294 => x"00011F6C",
000295 => x"00011F78",
000296 => x"00011F9C",
000297 => x"00011FA8",
000298 => x"00011FB4",
000299 => x"00011FB8",
000300 => x"00011FC8",
000301 => x"00011FDC",
000302 => x"E1A01000",
000303 => x"E5912000",
000304 => x"E59F0000",
000305 => x"EA000354",
000306 => x"00011FEC",
000307 => x"E2400001",
000308 => x"E92D4010",
000309 => x"E1A04001",
000310 => x"E3500004",
000311 => x"979FF100",
000312 => x"EA000039",
000313 => x"000104F8",
000314 => x"00010538",
000315 => x"0001054C",
000316 => x"00010578",
000317 => x"0001059C",
000318 => x"E59F10EC",
000319 => x"E59F00EC",
000320 => x"EB000345",
000321 => x"E3A01602",
000322 => x"E3A00505",
000323 => x"EB000153",
000324 => x"E3500602",
000325 => x"E1A04000",
000326 => x"81A01000",
000327 => x"8A000027",
000328 => x"E59F00CC",
000329 => x"EB00033C",
000330 => x"E1A01004",
000331 => x"E3A00505",
000332 => x"E8BD4010",
000333 => x"EA0001EE",
000334 => x"EBFFFF96",
000335 => x"EBFFFEDB",
000336 => x"E3A00010",
000337 => x"EBFFFF8A",
000338 => x"EA000008",
000339 => x"E3A01702",
000340 => x"E59F00A0",
000341 => x"EB000330",
000342 => x"E3A00010",
000343 => x"EBFFFF84",
000344 => x"E59F0094",
000345 => x"EB00032C",
000346 => x"E3A00702",
000347 => x"EBFFFEBD",
000348 => x"E8BD4010",
000349 => x"EA000346",
000350 => x"E3A01901",
000351 => x"E59F0074",
000352 => x"EB000325",
000353 => x"E3A00010",
000354 => x"EBFFFF79",
000355 => x"E59F0068",
000356 => x"EB000321",
000357 => x"E3A00901",
000358 => x"EAFFFFF3",
000359 => x"E59F1048",
000360 => x"E59F0048",
000361 => x"EB00031C",
000362 => x"E1A00004",
000363 => x"E3A01602",
000364 => x"EB00012A",
000365 => x"E3500602",
000366 => x"98BD8010",
000367 => x"E1A01000",
000368 => x"E59F0038",
000369 => x"E8BD4010",
000370 => x"EA000313",
000371 => x"E59F0024",
000372 => x"EB000311",
000373 => x"E3A00010",
000374 => x"EBFFFF65",
000375 => x"E59F0018",
000376 => x"EB00030D",
000377 => x"E1A00004",
000378 => x"EAFFFFDF",
000379 => x"00012008",
000380 => x"00012004",
000381 => x"00012068",
000382 => x"00012074",
000383 => x"00012064",
000384 => x"00012048",
000385 => x"E92D4010",
000386 => x"E59F3238",
000387 => x"E5D0C001",
000388 => x"E1A0E000",
000389 => x"E893000F",
000390 => x"E24DD020",
000391 => x"E35C0000",
000392 => x"E1A0400D",
000393 => x"E88D000F",
000394 => x"0A000084",
000395 => x"E35C000D",
000396 => x"1A000011",
000397 => x"E5DE0000",
000398 => x"E350006C",
000399 => x"0A000005",
000400 => x"E3500073",
000401 => x"0A000006",
000402 => x"E3500068",
000403 => x"1A00000C",
000404 => x"EBFFFF50",
000405 => x"EA000079",
000406 => x"E3A00001",
000407 => x"E3A01000",
000408 => x"EA000034",
000409 => x"EBFFFE91",
000410 => x"E3A00010",
000411 => x"EBFFFF40",
000412 => x"E59F01D4",
000413 => x"EB0002E8",
000414 => x"EA000070",
000415 => x"E35C0020",
000416 => x"0A000002",
000417 => x"E59F01C4",
000418 => x"E1A0100D",
000419 => x"EA00006A",
000420 => x"E5DE3000",
000421 => x"E353006A",
000422 => x"0A00001D",
000423 => x"8A000004",
000424 => x"E3530062",
000425 => x"0A00004D",
000426 => x"E3530064",
000427 => x"1A000060",
000428 => x"EA000006",
000429 => x"E3530072",
000430 => x"0A000040",
000431 => x"E3530077",
000432 => x"0A00004F",
000433 => x"E3530070",
000434 => x"1A000059",
000435 => x"EA00001B",
000436 => x"E1A0000E",
000437 => x"E28D1010",
000438 => x"E28D2014",
000439 => x"EBFFFF0F",
000440 => x"E3500000",
000441 => x"159D4010",
000442 => x"1A000001",
000443 => x"EA000053",
000444 => x"EBFFFF70",
000445 => x"E59D3010",
000446 => x"E59D2014",
000447 => x"E0833002",
000448 => x"E1540003",
000449 => x"E1A00004",
000450 => x"E2844004",
000451 => x"3AFFFFF7",
000452 => x"EA00004A",
000453 => x"E1A0000E",
000454 => x"E3A01002",
000455 => x"E28D2010",
000456 => x"E28D3018",
000457 => x"EBFFFE9E",
000458 => x"E3500000",
000459 => x"0A000043",
000460 => x"E3A00000",
000461 => x"E59D1010",
000462 => x"EBFFFF63",
000463 => x"EA00003F",
000464 => x"E1A0000E",
000465 => x"E3A01002",
000466 => x"E28D2010",
000467 => x"E28D3018",
000468 => x"EBFFFE93",
000469 => x"E3500000",
000470 => x"0A000038",
000471 => x"E3A03000",
000472 => x"E58D3018",
000473 => x"E59D3010",
000474 => x"E4D34001",
000475 => x"E58D3010",
000476 => x"EA00000B",
000477 => x"E3540000",
000478 => x"0A000003",
000479 => x"EB0002C8",
000480 => x"E354000D",
000481 => x"E59F00C0",
000482 => x"0B0002A3",
000483 => x"E59D2010",
000484 => x"E59D3018",
000485 => x"E4D24001",
000486 => x"E2833001",
000487 => x"E58D2010",
000488 => x"E58D3018",
000489 => x"E3140080",
000490 => x"E1A00004",
000491 => x"1A000023",
000492 => x"E59D3018",
000493 => x"E3530A01",
000494 => x"3AFFFFED",
000495 => x"EA00001F",
000496 => x"E1A0000E",
000497 => x"E3A01002",
000498 => x"E28D2010",
000499 => x"E28D3018",
000500 => x"EBFFFE73",
000501 => x"E3500000",
000502 => x"0A000018",
000503 => x"EA000011",
000504 => x"E1A0000E",
000505 => x"E3A01002",
000506 => x"E28D2010",
000507 => x"E28D3018",
000508 => x"EBFFFE6B",
000509 => x"E3500000",
000510 => x"13A00005",
000511 => x"1AFFFFCC",
000512 => x"EA00000E",
000513 => x"E1A0000E",
000514 => x"E28D1010",
000515 => x"E28D201C",
000516 => x"EBFFFEC2",
000517 => x"E3500000",
000518 => x"0A000008",
000519 => x"E59D201C",
000520 => x"E59D3010",
000521 => x"E5832000",
000522 => x"E59D0010",
000523 => x"EBFFFF21",
000524 => x"EA000002",
000525 => x"E59F0014",
000526 => x"E1A0100D",
000527 => x"EB000276",
000528 => x"E28DD020",
000529 => x"E8BD8010",
000530 => x"00012080",
000531 => x"00012064",
000532 => x"00012004",
000533 => x"E92D41F0",
000534 => x"E3A0100C",
000535 => x"E24DD028",
000536 => x"E59F2170",
000537 => x"E59F0170",
000538 => x"EB00026B",
000539 => x"EBFFFEC9",
000540 => x"E59F0168",
000541 => x"EB000268",
000542 => x"E3A06000",
000543 => x"E1A07006",
000544 => x"E1A08006",
000545 => x"EA000001",
000546 => x"E1A06008",
000547 => x"E3A07000",
000548 => x"E3A00FFA",
000549 => x"EB00028A",
000550 => x"E2504000",
000551 => x"BAFFFFFB",
000552 => x"E354001B",
000553 => x"0A00001C",
000554 => x"E3570001",
000555 => x"0354005B",
000556 => x"13A05000",
000557 => x"03A05001",
000558 => x"03A07002",
000559 => x"0A00001D",
000560 => x"E3570002",
000561 => x"1A000038",
000562 => x"E3540041",
000563 => x"01A04005",
000564 => x"11A07005",
000565 => x"1AFFFFED",
000566 => x"EA000000",
000567 => x"EB000270",
000568 => x"E1540006",
000569 => x"E3A00008",
000570 => x"E2844001",
000571 => x"BAFFFFFA",
000572 => x"E3A04000",
000573 => x"EA000005",
000574 => x"E28D3014",
000575 => x"E7D42003",
000576 => x"E1A00002",
000577 => x"E7C4200D",
000578 => x"EB000265",
000579 => x"E2844001",
000580 => x"E1540008",
000581 => x"BAFFFFF7",
000582 => x"EAFFFFDA",
000583 => x"E3A07001",
000584 => x"EA000004",
000585 => x"E28D2028",
000586 => x"E0823006",
000587 => x"E5434028",
000588 => x"E2866001",
000589 => x"E3A07000",
000590 => x"E3560012",
000591 => x"D3A03000",
000592 => x"C3A03001",
000593 => x"E354000D",
000594 => x"03833001",
000595 => x"E3530000",
000596 => x"0AFFFFCE",
000597 => x"E3560001",
000598 => x"DA000007",
000599 => x"E3A01000",
000600 => x"E7D1200D",
000601 => x"E28D3014",
000602 => x"E7C12003",
000603 => x"E2811001",
000604 => x"E3510014",
000605 => x"1AFFFFF9",
000606 => x"E2468001",
000607 => x"E28D2028",
000608 => x"E0823006",
000609 => x"E3A04000",
000610 => x"E5434028",
000611 => x"E59F0050",
000612 => x"EB000221",
000613 => x"E1A0000D",
000614 => x"EBFFFF19",
000615 => x"E59F0044",
000616 => x"EB00021D",
000617 => x"E1A06004",
000618 => x"EAFFFFB8",
000619 => x"EB00023C",
000620 => x"E3540008",
000621 => x"13A03000",
000622 => x"03A03001",
000623 => x"E3560000",
000624 => x"D3A03000",
000625 => x"E3530000",
000626 => x"12466001",
000627 => x"11A07005",
000628 => x"1AFFFFD8",
000629 => x"EAFFFFD2",
000630 => x"000120C4",
000631 => x"00012090",
000632 => x"000120D0",
000633 => x"00012064",
000634 => x"000120DC",
000635 => x"E92D4010",
000636 => x"E3A0C000",
000637 => x"E1A04000",
000638 => x"E1A0E00C",
000639 => x"E1A00001",
000640 => x"EA00000A",
000641 => x"E7DE3004",
000642 => x"E023342C",
000643 => x"E1A03083",
000644 => x"E0832001",
000645 => x"E7D31001",
000646 => x"E5D23001",
000647 => x"E1833401",
000648 => x"E023340C",
000649 => x"E1A03803",
000650 => x"E28EE001",
000651 => x"E1A0C823",
000652 => x"E15E0000",
000653 => x"E59F1008",
000654 => x"BAFFFFF1",
000655 => x"E1A0000C",
000656 => x"E8BD8010",
000657 => x"00011C44",
000658 => x"E52DE004",
000659 => x"E3A00F4B",
000660 => x"EB00021B",
000661 => x"E3500000",
000662 => x"AAFFFFFB",
000663 => x"E49DF004",
000664 => x"E92D4FF0",
000665 => x"E3A07000",
000666 => x"E24DDB01",
000667 => x"E24DD008",
000668 => x"E1A0B000",
000669 => x"E1A09001",
000670 => x"E3A0A019",
000671 => x"E3A04043",
000672 => x"E3A08001",
000673 => x"E1A06007",
000674 => x"EA000000",
000675 => x"E3A04015",
000676 => x"E3A05000",
000677 => x"E3540000",
000678 => x"11A00004",
000679 => x"1B000200",
000680 => x"E3A00FFA",
000681 => x"EB000206",
000682 => x"E3500000",
000683 => x"BA000019",
000684 => x"E3500002",
000685 => x"0A000025",
000686 => x"CA000002",
000687 => x"E3500001",
000688 => x"1A000014",
000689 => x"EA000004",
000690 => x"E3500004",
000691 => x"0A000004",
000692 => x"E3500018",
000693 => x"1A00000F",
000694 => x"EA000005",
000695 => x"E3A05080",
000696 => x"EA00001B",
000697 => x"E3A00006",
000698 => x"EB0001ED",
000699 => x"EBFFFFD5",
000700 => x"EA00007B",
000701 => x"E3A00FFA",
000702 => x"EB0001F1",
000703 => x"E3500018",
000704 => x"1A000004",
000705 => x"EBFFFFCF",
000706 => x"E3A00006",
000707 => x"EB0001E4",
000708 => x"E3E06000",
000709 => x"EA000072",
000710 => x"E2855001",
000711 => x"E3550050",
000712 => x"1AFFFFDB",
000713 => x"E3540043",
000714 => x"0AFFFFD7",
000715 => x"EBFFFFC5",
000716 => x"E3A00018",
000717 => x"EB0001DA",
000718 => x"E3A00018",
000719 => x"EB0001D8",
000720 => x"E3A00018",
000721 => x"EB0001D6",
000722 => x"E3E06001",
000723 => x"EA000064",
000724 => x"E3A05B01",
000725 => x"E3540043",
000726 => x"03A07001",
000727 => x"E1A00000",
000728 => x"E3A04000",
000729 => x"E5CD0002",
000730 => x"EA000006",
000731 => x"EB0001D4",
000732 => x"E28D3008",
000733 => x"E3500000",
000734 => x"E2433006",
000735 => x"E2844001",
000736 => x"BA000052",
000737 => x"E7C40003",
000738 => x"E3570000",
000739 => x"13A03004",
000740 => x"03A03003",
000741 => x"E0853003",
000742 => x"E1540003",
000743 => x"E3A00FFA",
000744 => x"BAFFFFF1",
000745 => x"E5DD3004",
000746 => x"E5DD2003",
000747 => x"E1E03003",
000748 => x"E20330FF",
000749 => x"E1520003",
000750 => x"1A000044",
000751 => x"E1520008",
000752 => x"0A000002",
000753 => x"E2483001",
000754 => x"E1520003",
000755 => x"1A00003F",
000756 => x"E3570000",
000757 => x"E28D4008",
000758 => x"E2444006",
000759 => x"01A01007",
000760 => x"02840003",
000761 => x"01A02001",
000762 => x"0A00000D",
000763 => x"E2840003",
000764 => x"E1A01005",
000765 => x"EBFFFF7C",
000766 => x"E0843005",
000767 => x"E5D32004",
000768 => x"E5D33003",
000769 => x"E0822403",
000770 => x"E1A02802",
000771 => x"E1500822",
000772 => x"1A00002E",
000773 => x"EA00000C",
000774 => x"E5503001",
000775 => x"E0813003",
000776 => x"E20310FF",
000777 => x"E1520005",
000778 => x"E2800001",
000779 => x"E2822001",
000780 => x"BAFFFFF8",
000781 => x"E28D2B01",
000782 => x"E2822008",
000783 => x"E0823005",
000784 => x"E5533403",
000785 => x"E1530001",
000786 => x"1A000020",
000787 => x"E5DD3003",
000788 => x"E1530008",
000789 => x"1A00000F",
000790 => x"E0663009",
000791 => x"E1550003",
000792 => x"B1A04005",
000793 => x"A1A04003",
000794 => x"E3540000",
000795 => x"DA000005",
000796 => x"E28D1008",
000797 => x"E08B0006",
000798 => x"E2411003",
000799 => x"E1A02004",
000800 => x"EB0002A0",
000801 => x"E0866004",
000802 => x"E2883001",
000803 => x"E20380FF",
000804 => x"E3A0A019",
000805 => x"EA00000B",
000806 => x"E24AA001",
000807 => x"E35A0000",
000808 => x"CA000008",
000809 => x"EBFFFF67",
000810 => x"E3A00018",
000811 => x"EB00017C",
000812 => x"E3A00018",
000813 => x"EB00017A",
000814 => x"E3A00018",
000815 => x"EB000178",
000816 => x"E3E06002",
000817 => x"EA000006",
000818 => x"E3A00006",
000819 => x"EA000001",
000820 => x"EBFFFF5C",
000821 => x"E3A00015",
000822 => x"EB000171",
000823 => x"E3A04000",
000824 => x"EAFFFF6A",
000825 => x"E1A00006",
000826 => x"E28DD008",
000827 => x"E28DDB01",
000828 => x"E8BD8FF0",
000829 => x"E92D40F0",
000830 => x"E59F1140",
000831 => x"E1A05000",
000832 => x"E3A02003",
000833 => x"E2800001",
000834 => x"EB00026A",
000835 => x"E3500000",
000836 => x"159F012C",
000837 => x"1A000006",
000838 => x"E5D52012",
000839 => x"E5D53013",
000840 => x"E1833402",
000841 => x"E3530028",
000842 => x"01A07000",
000843 => x"0A00003C",
000844 => x"E59F0110",
000845 => x"EB000138",
000846 => x"E3A00001",
000847 => x"E8BD80F0",
000848 => x"E5952020",
000849 => x"E5D5102E",
000850 => x"E5D5302F",
000851 => x"E0852002",
000852 => x"E1833401",
000853 => x"E0242397",
000854 => x"E5943004",
000855 => x"E3530001",
000856 => x"1A000018",
000857 => x"E5943014",
000858 => x"E3530000",
000859 => x"0A00002B",
000860 => x"E594300C",
000861 => x"E3530000",
000862 => x"13A06000",
000863 => x"1A00000E",
000864 => x"EA000026",
000865 => x"E5942010",
000866 => x"E0862002",
000867 => x"E0851002",
000868 => x"E5D13002",
000869 => x"E5D10003",
000870 => x"E7D5C002",
000871 => x"E1A03803",
000872 => x"E5D12001",
000873 => x"E1833C00",
000874 => x"E594E00C",
000875 => x"E183300C",
000876 => x"E1833402",
000877 => x"E78E3006",
000878 => x"E2866004",
000879 => x"E5943014",
000880 => x"E1560003",
000881 => x"3AFFFFEE",
000882 => x"E5943004",
000883 => x"E3530008",
000884 => x"1A000012",
000885 => x"E5943014",
000886 => x"E3530000",
000887 => x"0A00000F",
000888 => x"E594300C",
000889 => x"E3530000",
000890 => x"15941010",
000891 => x"1A000006",
000892 => x"EA00000A",
000893 => x"E594300C",
000894 => x"E0813003",
000895 => x"E0623003",
000896 => x"E3A02000",
000897 => x"E5832000",
000898 => x"E2811004",
000899 => x"E2842010",
000900 => x"E892000C",
000901 => x"E0823003",
000902 => x"E1510003",
000903 => x"3AFFFFF4",
000904 => x"E2877001",
000905 => x"E5D52030",
000906 => x"E5D53031",
000907 => x"E1833402",
000908 => x"E1570003",
000909 => x"3AFFFFC1",
000910 => x"E3A00000",
000911 => x"E8BD80F0",
000912 => x"000120E0",
000913 => x"000120E4",
000914 => x"00012100",
000915 => x"E5903000",
000916 => x"E20110FF",
000917 => x"E3530000",
000918 => x"14C31001",
000919 => x"E1A02000",
000920 => x"E1A00001",
000921 => x"15823000",
000922 => x"11A0F00E",
000923 => x"EA00010C",
000924 => x"E92D45F0",
000925 => x"E2525000",
000926 => x"E1A08000",
000927 => x"E1A07001",
000928 => x"C3A02000",
000929 => x"CA000001",
000930 => x"EA000009",
000931 => x"E2822001",
000932 => x"E7D21007",
000933 => x"E3510000",
000934 => x"1AFFFFFB",
000935 => x"E1520005",
000936 => x"A1A05001",
000937 => x"B0625005",
000938 => x"E3130002",
000939 => x"13A0A030",
000940 => x"1A000000",
000941 => x"E3A0A020",
000942 => x"E3130001",
000943 => x"13A06000",
000944 => x"01A04005",
000945 => x"0A000002",
000946 => x"EA00000A",
000947 => x"EBFFFFDE",
000948 => x"E2444001",
000949 => x"E3540000",
000950 => x"E1A00008",
000951 => x"E20A10FF",
000952 => x"CAFFFFF9",
000953 => x"E0646005",
000954 => x"E1A05004",
000955 => x"EA000001",
000956 => x"EBFFFFD5",
000957 => x"E2866001",
000958 => x"E5D73000",
000959 => x"E2531000",
000960 => x"E1A00008",
000961 => x"E2877001",
000962 => x"1AFFFFF8",
000963 => x"EA000001",
000964 => x"EBFFFFCD",
000965 => x"E2866001",
000966 => x"E3550000",
000967 => x"E1A00008",
000968 => x"E20A10FF",
000969 => x"E2455001",
000970 => x"CAFFFFF8",
000971 => x"E1A00006",
000972 => x"E8BD85F0",
000973 => x"E92D4FF0",
000974 => x"E2514000",
000975 => x"E24DD010",
000976 => x"E1A05002",
000977 => x"E1A09000",
000978 => x"E28D6034",
000979 => x"E8960C40",
000980 => x"1A000007",
000981 => x"E3A0C030",
000982 => x"E1A02006",
000983 => x"E1A0300A",
000984 => x"E1A0100D",
000985 => x"E5CDC000",
000986 => x"E5CD4001",
000987 => x"EBFFFFBF",
000988 => x"EA00003C",
000989 => x"E2533000",
000990 => x"13A03001",
000991 => x"E352000A",
000992 => x"13A03000",
000993 => x"E3530000",
000994 => x"0A000003",
000995 => x"E3540000",
000996 => x"B2644000",
000997 => x"B3A08001",
000998 => x"BA000000",
000999 => x"E3A08000",
001000 => x"E3A03000",
001001 => x"E28D700F",
001002 => x"E5CD300F",
001003 => x"EA000010",
001004 => x"E3550010",
001005 => x"0A000002",
001006 => x"EB0000CD",
001007 => x"E0030095",
001008 => x"E0633004",
001009 => x"E3530009",
001010 => x"E083200B",
001011 => x"C242303A",
001012 => x"E2833030",
001013 => x"E3550010",
001014 => x"E1A00004",
001015 => x"E1A01005",
001016 => x"E5673001",
001017 => x"01A04224",
001018 => x"0A000001",
001019 => x"EB0000C0",
001020 => x"E1A04000",
001021 => x"E3540000",
001022 => x"E1A00004",
001023 => x"E1A01005",
001024 => x"E204300F",
001025 => x"1AFFFFE9",
001026 => x"E3580000",
001027 => x"E1A02007",
001028 => x"01A04008",
001029 => x"0A00000D",
001030 => x"E3560000",
001031 => x"0A000007",
001032 => x"E31A0002",
001033 => x"0A000005",
001034 => x"E1A00009",
001035 => x"E3A0102D",
001036 => x"EBFFFF85",
001037 => x"E2466001",
001038 => x"E3A04001",
001039 => x"EA000003",
001040 => x"E3A0302D",
001041 => x"E5423001",
001042 => x"E2477001",
001043 => x"E3A04000",
001044 => x"E1A00009",
001045 => x"E1A01007",
001046 => x"E1A02006",
001047 => x"E1A0300A",
001048 => x"EBFFFF82",
001049 => x"E0840000",
001050 => x"E28DD010",
001051 => x"E8BD8FF0",
001052 => x"E92D41F0",
001053 => x"E1A07000",
001054 => x"E24DD010",
001055 => x"E1A04001",
001056 => x"E1A05002",
001057 => x"E3A06000",
001058 => x"EA00005C",
001059 => x"E3530025",
001060 => x"1A000051",
001061 => x"E5F43001",
001062 => x"E3530000",
001063 => x"0A00005A",
001064 => x"E3530025",
001065 => x"0A000050",
001066 => x"E353002D",
001067 => x"13A08000",
001068 => x"02844001",
001069 => x"03A08001",
001070 => x"EA000001",
001071 => x"E2844001",
001072 => x"E3888002",
001073 => x"E5D43000",
001074 => x"E3530030",
001075 => x"0AFFFFFA",
001076 => x"E3A0E000",
001077 => x"EA000003",
001078 => x"E3A0300A",
001079 => x"E023239E",
001080 => x"E2844001",
001081 => x"E243E030",
001082 => x"E5D42000",
001083 => x"E2423030",
001084 => x"E3530009",
001085 => x"9AFFFFF7",
001086 => x"E3520073",
001087 => x"1A000007",
001088 => x"E4953004",
001089 => x"E59F110C",
001090 => x"E3530000",
001091 => x"11A01003",
001092 => x"E1A0200E",
001093 => x"E1A03008",
001094 => x"E1A00007",
001095 => x"EA00002C",
001096 => x"E3520064",
001097 => x"1A00000A",
001098 => x"E4951004",
001099 => x"E1A00007",
001100 => x"E3A0200A",
001101 => x"E3A03001",
001102 => x"E58DE000",
001103 => x"E58D8004",
001104 => x"E3A0C061",
001105 => x"E58DC008",
001106 => x"EBFFFF79",
001107 => x"E0866000",
001108 => x"EA000029",
001109 => x"E3520078",
001110 => x"04951004",
001111 => x"01A00007",
001112 => x"03A02010",
001113 => x"0A00000E",
001114 => x"E3520058",
001115 => x"1A000007",
001116 => x"E4951004",
001117 => x"E1A00007",
001118 => x"E3A02010",
001119 => x"E3A03000",
001120 => x"E3A0C041",
001121 => x"E58DE000",
001122 => x"E58D8004",
001123 => x"EAFFFFEC",
001124 => x"E3520075",
001125 => x"1A000004",
001126 => x"E4951004",
001127 => x"E1A00007",
001128 => x"E3A0200A",
001129 => x"E3A03000",
001130 => x"EAFFFFE2",
001131 => x"E3520063",
001132 => x"1A000011",
001133 => x"E495C004",
001134 => x"E5CDC00E",
001135 => x"E3A0C000",
001136 => x"E5CDC00F",
001137 => x"E1A0200E",
001138 => x"E1A03008",
001139 => x"E1A00007",
001140 => x"E28D100E",
001141 => x"EBFFFF25",
001142 => x"EAFFFFDB",
001143 => x"E353000A",
001144 => x"01A00007",
001145 => x"03A0100D",
001146 => x"0BFFFF17",
001147 => x"E1A00007",
001148 => x"E5D41000",
001149 => x"EBFFFF14",
001150 => x"E2866001",
001151 => x"E2844001",
001152 => x"E5D43000",
001153 => x"E3530000",
001154 => x"1AFFFF9F",
001155 => x"E1A00006",
001156 => x"E28DD010",
001157 => x"E8BD81F0",
001158 => x"00012138",
001159 => x"E92D000F",
001160 => x"E52DE004",
001161 => x"E24DD004",
001162 => x"E28D0004",
001163 => x"E3A03000",
001164 => x"E5203004",
001165 => x"E59D1008",
001166 => x"E1A0000D",
001167 => x"E28D200C",
001168 => x"EBFFFF8A",
001169 => x"E28DD004",
001170 => x"E49DE004",
001171 => x"E28DD010",
001172 => x"E1A0F00E",
001173 => x"E92D000E",
001174 => x"E52DE004",
001175 => x"E24DD004",
001176 => x"E28D3004",
001177 => x"E5230004",
001178 => x"E59D1008",
001179 => x"E1A0000D",
001180 => x"E28D200C",
001181 => x"EBFFFF7D",
001182 => x"E28DD004",
001183 => x"E49DE004",
001184 => x"E28DD00C",
001185 => x"E1A0F00E",
001186 => x"E59FB46C",
001187 => x"E58B0000",
001188 => x"EAFFFFFC",
001189 => x"E59FB460",
001190 => x"E3A0A011",
001191 => x"E58BA000",
001192 => x"EAFFFFFB",
001193 => x"E59F1454",
001194 => x"E59F3454",
001195 => x"E5932000",
001196 => x"E2022020",
001197 => x"E3520000",
001198 => x"05810000",
001199 => x"01B0F00E",
001200 => x"1AFFFFF9",
001201 => x"E59F2434",
001202 => x"E59F3434",
001203 => x"E1A01580",
001204 => x"E0811480",
001205 => x"E5930000",
001206 => x"E2100010",
001207 => x"05920000",
001208 => x"01A0F00E",
001209 => x"E2511001",
001210 => x"1AFFFFF9",
001211 => x"E3E00000",
001212 => x"E1B0F00E",
001213 => x"E92D4010",
001214 => x"E2002102",
001215 => x"E2013102",
001216 => x"E0224003",
001217 => x"E3100102",
001218 => x"11E00000",
001219 => x"12800001",
001220 => x"E3110102",
001221 => x"11E01001",
001222 => x"12811001",
001223 => x"E1A02001",
001224 => x"E1A01000",
001225 => x"E3520000",
001226 => x"0A000011",
001227 => x"E3A00000",
001228 => x"E3A03001",
001229 => x"E3530000",
001230 => x"03A03201",
001231 => x"0A000003",
001232 => x"E1520001",
001233 => x"91A02082",
001234 => x"91A03083",
001235 => x"9AFFFFF8",
001236 => x"E1510002",
001237 => x"20411002",
001238 => x"20800003",
001239 => x"E1B030A3",
001240 => x"31A020A2",
001241 => x"3AFFFFF9",
001242 => x"E3140102",
001243 => x"11E00000",
001244 => x"12800001",
001245 => x"E8FD8010",
001246 => x"E92D4070",
001247 => x"E1A06000",
001248 => x"E1862001",
001249 => x"E3120003",
001250 => x"1A00002A",
001251 => x"E8B1003C",
001252 => x"E31200FF",
001253 => x"13120CFF",
001254 => x"131208FF",
001255 => x"131204FF",
001256 => x"14862004",
001257 => x"02411004",
001258 => x"131300FF",
001259 => x"13130CFF",
001260 => x"131308FF",
001261 => x"131304FF",
001262 => x"14863004",
001263 => x"02411004",
001264 => x"131400FF",
001265 => x"13140CFF",
001266 => x"131408FF",
001267 => x"131404FF",
001268 => x"14864004",
001269 => x"02411004",
001270 => x"131500FF",
001271 => x"13150CFF",
001272 => x"131508FF",
001273 => x"131504FF",
001274 => x"14865004",
001275 => x"02411004",
001276 => x"1AFFFFE5",
001277 => x"E4913004",
001278 => x"E4C63001",
001279 => x"E21340FF",
001280 => x"08FD8070",
001281 => x"E1A03423",
001282 => x"E4C63001",
001283 => x"E21340FF",
001284 => x"08FD8070",
001285 => x"E1A03423",
001286 => x"E4C63001",
001287 => x"E21340FF",
001288 => x"08FD8070",
001289 => x"E1A03423",
001290 => x"E4C63001",
001291 => x"E21340FF",
001292 => x"08FD8070",
001293 => x"EAFFFFEE",
001294 => x"E4D13001",
001295 => x"E4C63001",
001296 => x"E3530000",
001297 => x"08FD8070",
001298 => x"E4D13001",
001299 => x"E4C63001",
001300 => x"E3530000",
001301 => x"08FD8070",
001302 => x"E4D13001",
001303 => x"E4C63001",
001304 => x"E3530000",
001305 => x"08FD8070",
001306 => x"E4D13001",
001307 => x"E4C63001",
001308 => x"E3530000",
001309 => x"08FD8070",
001310 => x"EAFFFFEE",
001311 => x"E92D41F0",
001312 => x"E1802001",
001313 => x"E3120003",
001314 => x"1A000018",
001315 => x"E8B0001C",
001316 => x"E8B100E0",
001317 => x"E1520005",
001318 => x"1A000012",
001319 => x"01530006",
001320 => x"1A00002B",
001321 => x"01540007",
001322 => x"1A000049",
001323 => x"E31200FF",
001324 => x"13120CFF",
001325 => x"131208FF",
001326 => x"131204FF",
001327 => x"131300FF",
001328 => x"13130CFF",
001329 => x"131308FF",
001330 => x"131304FF",
001331 => x"131400FF",
001332 => x"13140CFF",
001333 => x"131408FF",
001334 => x"131404FF",
001335 => x"1AFFFFEA",
001336 => x"03A00000",
001337 => x"08FD81F0",
001338 => x"E240000C",
001339 => x"E241100C",
001340 => x"E4D02001",
001341 => x"E4D13001",
001342 => x"E0324003",
001343 => x"1A00005A",
001344 => x"E4D05001",
001345 => x"E4D16001",
001346 => x"E3520000",
001347 => x"0A000054",
001348 => x"E0357006",
001349 => x"1A000054",
001350 => x"E4D02001",
001351 => x"E4D13001",
001352 => x"E3550000",
001353 => x"0A00004E",
001354 => x"E0324003",
001355 => x"1A00004E",
001356 => x"E4D05001",
001357 => x"E4D16001",
001358 => x"E3520000",
001359 => x"0A000048",
001360 => x"E0357006",
001361 => x"1A000048",
001362 => x"E3550000",
001363 => x"0A000044",
001364 => x"1AFFFFE6",
001365 => x"E31200FF",
001366 => x"13120CFF",
001367 => x"131208FF",
001368 => x"131204FF",
001369 => x"0A00003E",
001370 => x"E2400008",
001371 => x"E2411008",
001372 => x"E4D02001",
001373 => x"E4D13001",
001374 => x"E0324003",
001375 => x"1A00003A",
001376 => x"E4D05001",
001377 => x"E4D16001",
001378 => x"E3520000",
001379 => x"0A000034",
001380 => x"E0357006",
001381 => x"1A000034",
001382 => x"E4D02001",
001383 => x"E4D13001",
001384 => x"E3550000",
001385 => x"0A00002E",
001386 => x"E0324003",
001387 => x"1A00002E",
001388 => x"E4D05001",
001389 => x"E4D16001",
001390 => x"E3520000",
001391 => x"0A000028",
001392 => x"E0357006",
001393 => x"1A000028",
001394 => x"E3550000",
001395 => x"0A000024",
001396 => x"1AFFFFC6",
001397 => x"E31200FF",
001398 => x"13120CFF",
001399 => x"131208FF",
001400 => x"131204FF",
001401 => x"131300FF",
001402 => x"13130CFF",
001403 => x"131308FF",
001404 => x"131304FF",
001405 => x"0A00001A",
001406 => x"E2400004",
001407 => x"E2411004",
001408 => x"E4D02001",
001409 => x"E4D13001",
001410 => x"E0324003",
001411 => x"1A000016",
001412 => x"E4D05001",
001413 => x"E4D16001",
001414 => x"E3520000",
001415 => x"0A000010",
001416 => x"E0357006",
001417 => x"1A000010",
001418 => x"E4D02001",
001419 => x"E4D13001",
001420 => x"E3550000",
001421 => x"0A00000A",
001422 => x"E0324003",
001423 => x"1A00000A",
001424 => x"E4D05001",
001425 => x"E4D16001",
001426 => x"E3520000",
001427 => x"0A000004",
001428 => x"E0357006",
001429 => x"1A000004",
001430 => x"E3550000",
001431 => x"0A000000",
001432 => x"1AFFFFA2",
001433 => x"03A00000",
001434 => x"08FD81F0",
001435 => x"E0450006",
001436 => x"E8FD81F0",
001437 => x"E59F107C",
001438 => x"E5811000",
001439 => x"E1A0F00E",
001440 => x"E59F1070",
001441 => x"E5910000",
001442 => x"E2800801",
001443 => x"E5810000",
001444 => x"E1A0F00E",
001445 => x"E92D4010",
001446 => x"E3520000",
001447 => x"0A000004",
001448 => x"E0804002",
001449 => x"E4D13001",
001450 => x"E4C03001",
001451 => x"E1500004",
001452 => x"1AFFFFFB",
001453 => x"E8FD8010",
001454 => x"E92D4070",
001455 => x"E3520000",
001456 => x"03A00001",
001457 => x"0A00000A",
001458 => x"E3A03000",
001459 => x"E2833001",
001460 => x"E4D04001",
001461 => x"E4D15001",
001462 => x"E0546005",
001463 => x"11A00006",
001464 => x"1A000003",
001465 => x"E1530002",
001466 => x"03A00000",
001467 => x"0A000000",
001468 => x"EAFFFFF5",
001469 => x"E8FD8070",
001470 => x"07000000",
001471 => x"F0000000",
001472 => x"FFFF0200",
001473 => x"FFFF0218",
001474 => x"E3520007",
001475 => x"E92D45F0",
001476 => x"E1A0C001",
001477 => x"E1A04002",
001478 => x"E1A0A000",
001479 => x"E1A0E000",
001480 => x"83A02000",
001481 => x"8A00001E",
001482 => x"E2443001",
001483 => x"E3530006",
001484 => x"979FF103",
001485 => x"EA000140",
001486 => x"0001178C",
001487 => x"00011784",
001488 => x"0001177C",
001489 => x"00011774",
001490 => x"0001176C",
001491 => x"00011764",
001492 => x"00011754",
001493 => x"E4D13001",
001494 => x"E1A0E000",
001495 => x"E4CE3001",
001496 => x"E1A0C001",
001497 => x"E4DC3001",
001498 => x"E4CE3001",
001499 => x"E4DC3001",
001500 => x"E4CE3001",
001501 => x"E4DC3001",
001502 => x"E4CE3001",
001503 => x"E4DC3001",
001504 => x"E4CE3001",
001505 => x"E4DC3001",
001506 => x"E4CE3001",
001507 => x"E5DC3000",
001508 => x"E5CE3000",
001509 => x"EA000128",
001510 => x"E7D23001",
001511 => x"E7C2300A",
001512 => x"E2822001",
001513 => x"E08AE002",
001514 => x"E31E0003",
001515 => x"1AFFFFF9",
001516 => x"E0811002",
001517 => x"E2013003",
001518 => x"E0626004",
001519 => x"E3530003",
001520 => x"979FF103",
001521 => x"EA00011B",
001522 => x"000117D8",
001523 => x"000118A8",
001524 => x"000119B8",
001525 => x"00011AC8",
001526 => x"E1A02126",
001527 => x"E3A0C000",
001528 => x"EA000003",
001529 => x"E79C3001",
001530 => x"E2422001",
001531 => x"E78C300E",
001532 => x"E28CC004",
001533 => x"E3120007",
001534 => x"1AFFFFF9",
001535 => x"E08E500C",
001536 => x"E081100C",
001537 => x"E1A021A2",
001538 => x"E1A0E005",
001539 => x"E1A0C001",
001540 => x"E1A04002",
001541 => x"EA00000F",
001542 => x"E51C3020",
001543 => x"E50E3020",
001544 => x"E51C301C",
001545 => x"E50E301C",
001546 => x"E51C3018",
001547 => x"E50E3018",
001548 => x"E51C3014",
001549 => x"E50E3014",
001550 => x"E51C3010",
001551 => x"E50E3010",
001552 => x"E51C300C",
001553 => x"E50E300C",
001554 => x"E51C3008",
001555 => x"E50E3008",
001556 => x"E51C3004",
001557 => x"E50E3004",
001558 => x"E2444001",
001559 => x"E3740001",
001560 => x"E28EE020",
001561 => x"E28CC020",
001562 => x"1AFFFFEA",
001563 => x"E2063003",
001564 => x"E1A02282",
001565 => x"E2433001",
001566 => x"E085C002",
001567 => x"E0811002",
001568 => x"E3530006",
001569 => x"979FF103",
001570 => x"EA0000EB",
001571 => x"00011C2C",
001572 => x"00011C24",
001573 => x"00011C1C",
001574 => x"00011C14",
001575 => x"00011C0C",
001576 => x"00011C04",
001577 => x"00011BFC",
001578 => x"E3C10003",
001579 => x"E5904000",
001580 => x"E3CE1003",
001581 => x"E1A0C126",
001582 => x"E1A02001",
001583 => x"EA000003",
001584 => x"E7954003",
001585 => x"E18E3C04",
001586 => x"E5023004",
001587 => x"E24CC001",
001588 => x"E2822004",
001589 => x"E31C0007",
001590 => x"E2615000",
001591 => x"E1A0E424",
001592 => x"E0803002",
001593 => x"1AFFFFF5",
001594 => x"E0613000",
001595 => x"E0837002",
001596 => x"E1A001AC",
001597 => x"E2428004",
001598 => x"E1A0E008",
001599 => x"E1A0C007",
001600 => x"E1A05000",
001601 => x"EA00001F",
001602 => x"E51C2020",
001603 => x"E1A03C02",
001604 => x"E1833424",
001605 => x"E50E3020",
001606 => x"E51C101C",
001607 => x"E1A03C01",
001608 => x"E1833422",
001609 => x"E50E301C",
001610 => x"E51C2018",
001611 => x"E1A03C02",
001612 => x"E1833421",
001613 => x"E50E3018",
001614 => x"E51C1014",
001615 => x"E1A03C01",
001616 => x"E1833422",
001617 => x"E50E3014",
001618 => x"E51C2010",
001619 => x"E1A03C02",
001620 => x"E1833421",
001621 => x"E50E3010",
001622 => x"E51C100C",
001623 => x"E1A03C01",
001624 => x"E1833422",
001625 => x"E50E300C",
001626 => x"E51C2008",
001627 => x"E1A03C02",
001628 => x"E1833421",
001629 => x"E50E3008",
001630 => x"E51C4004",
001631 => x"E1A03C04",
001632 => x"E1833422",
001633 => x"E50E3004",
001634 => x"E2455001",
001635 => x"E3750001",
001636 => x"E28EE020",
001637 => x"E28CC020",
001638 => x"1AFFFFDA",
001639 => x"E1A03280",
001640 => x"E2062003",
001641 => x"E0871003",
001642 => x"E2422001",
001643 => x"E088C003",
001644 => x"E2411003",
001645 => x"EA000086",
001646 => x"E3C10003",
001647 => x"E5904000",
001648 => x"E3CE1003",
001649 => x"E1A0C126",
001650 => x"E1A02001",
001651 => x"EA000003",
001652 => x"E7954003",
001653 => x"E18E3804",
001654 => x"E5023004",
001655 => x"E24CC001",
001656 => x"E2822004",
001657 => x"E31C0007",
001658 => x"E2615000",
001659 => x"E1A0E824",
001660 => x"E0803002",
001661 => x"1AFFFFF5",
001662 => x"E0613000",
001663 => x"E0837002",
001664 => x"E1A001AC",
001665 => x"E2428004",
001666 => x"E1A0E008",
001667 => x"E1A0C007",
001668 => x"E1A05000",
001669 => x"EA00001F",
001670 => x"E51C2020",
001671 => x"E1A03802",
001672 => x"E1833824",
001673 => x"E50E3020",
001674 => x"E51C101C",
001675 => x"E1A03801",
001676 => x"E1833822",
001677 => x"E50E301C",
001678 => x"E51C2018",
001679 => x"E1A03802",
001680 => x"E1833821",
001681 => x"E50E3018",
001682 => x"E51C1014",
001683 => x"E1A03801",
001684 => x"E1833822",
001685 => x"E50E3014",
001686 => x"E51C2010",
001687 => x"E1A03802",
001688 => x"E1833821",
001689 => x"E50E3010",
001690 => x"E51C100C",
001691 => x"E1A03801",
001692 => x"E1833822",
001693 => x"E50E300C",
001694 => x"E51C2008",
001695 => x"E1A03802",
001696 => x"E1833821",
001697 => x"E50E3008",
001698 => x"E51C4004",
001699 => x"E1A03804",
001700 => x"E1833822",
001701 => x"E50E3004",
001702 => x"E2455001",
001703 => x"E3750001",
001704 => x"E28EE020",
001705 => x"E28CC020",
001706 => x"1AFFFFDA",
001707 => x"E1A03280",
001708 => x"E2062003",
001709 => x"E0871003",
001710 => x"E2422001",
001711 => x"E088C003",
001712 => x"E2411002",
001713 => x"EA000042",
001714 => x"E3C10003",
001715 => x"E5904000",
001716 => x"E3CE1003",
001717 => x"E1A0C126",
001718 => x"E1A02001",
001719 => x"EA000003",
001720 => x"E7954003",
001721 => x"E18E3404",
001722 => x"E5023004",
001723 => x"E24CC001",
001724 => x"E2822004",
001725 => x"E31C0007",
001726 => x"E2615000",
001727 => x"E1A0EC24",
001728 => x"E0803002",
001729 => x"1AFFFFF5",
001730 => x"E0613000",
001731 => x"E0837002",
001732 => x"E1A001AC",
001733 => x"E2428004",
001734 => x"E1A0E008",
001735 => x"E1A0C007",
001736 => x"E1A05000",
001737 => x"EA00001F",
001738 => x"E51C2020",
001739 => x"E1A03402",
001740 => x"E1833C24",
001741 => x"E50E3020",
001742 => x"E51C101C",
001743 => x"E1A03401",
001744 => x"E1833C22",
001745 => x"E50E301C",
001746 => x"E51C2018",
001747 => x"E1A03402",
001748 => x"E1833C21",
001749 => x"E50E3018",
001750 => x"E51C1014",
001751 => x"E1A03401",
001752 => x"E1833C22",
001753 => x"E50E3014",
001754 => x"E51C2010",
001755 => x"E1A03402",
001756 => x"E1833C21",
001757 => x"E50E3010",
001758 => x"E51C100C",
001759 => x"E1A03401",
001760 => x"E1833C22",
001761 => x"E50E300C",
001762 => x"E51C2008",
001763 => x"E1A03402",
001764 => x"E1833C21",
001765 => x"E50E3008",
001766 => x"E51C4004",
001767 => x"E1A03404",
001768 => x"E1833C22",
001769 => x"E50E3004",
001770 => x"E2455001",
001771 => x"E3750001",
001772 => x"E28EE020",
001773 => x"E28CC020",
001774 => x"1AFFFFDA",
001775 => x"E1A03280",
001776 => x"E2062003",
001777 => x"E0871003",
001778 => x"E2422001",
001779 => x"E088C003",
001780 => x"E2411001",
001781 => x"E3520006",
001782 => x"979FF102",
001783 => x"EA000016",
001784 => x"00011C2C",
001785 => x"00011C24",
001786 => x"00011C1C",
001787 => x"00011C14",
001788 => x"00011C0C",
001789 => x"00011C04",
001790 => x"00011BFC",
001791 => x"E4D13001",
001792 => x"E4CC3001",
001793 => x"E4D13001",
001794 => x"E4CC3001",
001795 => x"E4D13001",
001796 => x"E4CC3001",
001797 => x"E4D13001",
001798 => x"E4CC3001",
001799 => x"E4D13001",
001800 => x"E4CC3001",
001801 => x"E4D13001",
001802 => x"E4CC3001",
001803 => x"E5D13000",
001804 => x"E5CC3000",
001805 => x"EA000000",
001806 => x"E8BD85F0",
001807 => x"E1A0000A",
001808 => x"E8BD85F0",
001809 => x"00001021",
001810 => x"20423063",
001811 => x"408450A5",
001812 => x"60C670E7",
001813 => x"81089129",
001814 => x"A14AB16B",
001815 => x"C18CD1AD",
001816 => x"E1CEF1EF",
001817 => x"12310210",
001818 => x"32732252",
001819 => x"52B54294",
001820 => x"72F762D6",
001821 => x"93398318",
001822 => x"B37BA35A",
001823 => x"D3BDC39C",
001824 => x"F3FFE3DE",
001825 => x"24623443",
001826 => x"04201401",
001827 => x"64E674C7",
001828 => x"44A45485",
001829 => x"A56AB54B",
001830 => x"85289509",
001831 => x"E5EEF5CF",
001832 => x"C5ACD58D",
001833 => x"36532672",
001834 => x"16110630",
001835 => x"76D766F6",
001836 => x"569546B4",
001837 => x"B75BA77A",
001838 => x"97198738",
001839 => x"F7DFE7FE",
001840 => x"D79DC7BC",
001841 => x"48C458E5",
001842 => x"688678A7",
001843 => x"08401861",
001844 => x"28023823",
001845 => x"C9CCD9ED",
001846 => x"E98EF9AF",
001847 => x"89489969",
001848 => x"A90AB92B",
001849 => x"5AF54AD4",
001850 => x"7AB76A96",
001851 => x"1A710A50",
001852 => x"3A332A12",
001853 => x"DBFDCBDC",
001854 => x"FBBFEB9E",
001855 => x"9B798B58",
001856 => x"BB3BAB1A",
001857 => x"6CA67C87",
001858 => x"4CE45CC5",
001859 => x"2C223C03",
001860 => x"0C601C41",
001861 => x"EDAEFD8F",
001862 => x"CDECDDCD",
001863 => x"AD2ABD0B",
001864 => x"8D689D49",
001865 => x"7E976EB6",
001866 => x"5ED54EF4",
001867 => x"3E132E32",
001868 => x"1E510E70",
001869 => x"FF9FEFBE",
001870 => x"DFDDCFFC",
001871 => x"BF1BAF3A",
001872 => x"9F598F78",
001873 => x"918881A9",
001874 => x"B1CAA1EB",
001875 => x"D10CC12D",
001876 => x"F14EE16F",
001877 => x"108000A1",
001878 => x"30C220E3",
001879 => x"50044025",
001880 => x"70466067",
001881 => x"83B99398",
001882 => x"A3FBB3DA",
001883 => x"C33DD31C",
001884 => x"E37FF35E",
001885 => x"02B11290",
001886 => x"22F332D2",
001887 => x"42355214",
001888 => x"62777256",
001889 => x"B5EAA5CB",
001890 => x"95A88589",
001891 => x"F56EE54F",
001892 => x"D52CC50D",
001893 => x"34E224C3",
001894 => x"14A00481",
001895 => x"74666447",
001896 => x"54244405",
001897 => x"A7DBB7FA",
001898 => x"879997B8",
001899 => x"E75FF77E",
001900 => x"C71DD73C",
001901 => x"26D336F2",
001902 => x"069116B0",
001903 => x"66577676",
001904 => x"46155634",
001905 => x"D94CC96D",
001906 => x"F90EE92F",
001907 => x"99C889E9",
001908 => x"B98AA9AB",
001909 => x"58444865",
001910 => x"78066827",
001911 => x"18C008E1",
001912 => x"388228A3",
001913 => x"CB7DDB5C",
001914 => x"EB3FFB1E",
001915 => x"8BF99BD8",
001916 => x"ABBBBB9A",
001917 => x"4A755A54",
001918 => x"6A377A16",
001919 => x"0AF11AD0",
001920 => x"2AB33A92",
001921 => x"FD2EED0F",
001922 => x"DD6CCD4D",
001923 => x"BDAAAD8B",
001924 => x"9DE88DC9",
001925 => x"7C266C07",
001926 => x"5C644C45",
001927 => x"3CA22C83",
001928 => x"1CE00CC1",
001929 => x"EF1FFF3E",
001930 => x"CF5DDF7C",
001931 => x"AF9BBFBA",
001932 => x"8FD99FF8",
001933 => x"6E177E36",
001934 => x"4E555E74",
001935 => x"2E933EB2",
001936 => x"0ED11EF0",
001937 => x"2573200A",
001938 => x"00000000",
001939 => x"63686172",
001940 => x"3A202563",
001941 => x"20000000",
001942 => x"30207468",
001943 => x"72752039",
001944 => x"00000000",
001945 => x"41207468",
001946 => x"72752046",
001947 => x"00000000",
001948 => x"61207468",
001949 => x"72752066",
001950 => x"00000000",
001951 => x"63706F73",
001952 => x"3A257820",
001953 => x"00000000",
001954 => x"61646472",
001955 => x"3A25780A",
001956 => x"00000000",
001957 => x"25692000",
001958 => x"436F6D6D",
001959 => x"616E6473",
001960 => x"0A000000",
001961 => x"6C000000",
001962 => x"3A204C6F",
001963 => x"61642065",
001964 => x"6C662066",
001965 => x"696C650A",
001966 => x"00000000",
001967 => x"62203C61",
001968 => x"64647265",
001969 => x"73733E00",
001970 => x"3A204C6F",
001971 => x"61642062",
001972 => x"696E6172",
001973 => x"79206669",
001974 => x"6C652074",
001975 => x"6F203C61",
001976 => x"64647265",
001977 => x"73733E0A",
001978 => x"00000000",
001979 => x"64203C73",
001980 => x"74617274",
001981 => x"20616464",
001982 => x"72657373",
001983 => x"3E203C6E",
001984 => x"756D2062",
001985 => x"79746573",
001986 => x"3E203A20",
001987 => x"44756D70",
001988 => x"206D656D",
001989 => x"0A000000",
001990 => x"68000000",
001991 => x"3A205072",
001992 => x"696E7420",
001993 => x"68656C70",
001994 => x"206D6573",
001995 => x"73616765",
001996 => x"0A000000",
001997 => x"6A203C61",
001998 => x"64647265",
001999 => x"73733E00",
002000 => x"3A204578",
002001 => x"65637574",
002002 => x"65206C6F",
002003 => x"61646564",
002004 => x"20656C66",
002005 => x"2C206A75",
002006 => x"6D70696E",
002007 => x"6720746F",
002008 => x"203C6164",
002009 => x"64726573",
002010 => x"733E0A00",
002011 => x"70203C61",
002012 => x"64647265",
002013 => x"73733E00",
002014 => x"3A205072",
002015 => x"696E7420",
002016 => x"61736369",
002017 => x"69206D65",
002018 => x"6D20756E",
002019 => x"74696C20",
002020 => x"66697273",
002021 => x"7420300A",
002022 => x"00000000",
002023 => x"72203C61",
002024 => x"64647265",
002025 => x"73733E00",
002026 => x"3A205265",
002027 => x"6164206D",
002028 => x"656D0A00",
002029 => x"73000000",
002030 => x"3A20436F",
002031 => x"72652073",
002032 => x"74617475",
002033 => x"730A0000",
002034 => x"77203C61",
002035 => x"64647265",
002036 => x"73733E20",
002037 => x"3C76616C",
002038 => x"75653E00",
002039 => x"3A205772",
002040 => x"69746520",
002041 => x"6D656D0A",
002042 => x"00000000",
002043 => x"6D656D20",
002044 => x"30782530",
002045 => x"3878203D",
002046 => x"20307825",
002047 => x"3038780A",
002048 => x"00000000",
002049 => x"25730A00",
002050 => x"53656E64",
002051 => x"2066696C",
002052 => x"6520772F",
002053 => x"20314B20",
002054 => x"586D6F64",
002055 => x"656D2070",
002056 => x"726F746F",
002057 => x"636F6C20",
002058 => x"66726F6D",
002059 => x"20746572",
002060 => x"6D696E61",
002061 => x"6C20656D",
002062 => x"756C6174",
002063 => x"6F72206E",
002064 => x"6F772E2E",
002065 => x"2E000000",
002066 => x"586D6F64",
002067 => x"656D2065",
002068 => x"72726F72",
002069 => x"2066696C",
002070 => x"65207369",
002071 => x"7A652030",
002072 => x"78257820",
002073 => x"0A000000",
002074 => x"0A656C66",
002075 => x"2073706C",
002076 => x"69740A00",
002077 => x"6A203078",
002078 => x"25303878",
002079 => x"0A000000",
002080 => x"496E7661",
002081 => x"6C696420",
002082 => x"636F6D6D",
002083 => x"616E6400",
002084 => x"2563416D",
002085 => x"62657220",
002086 => x"426F6F74",
002087 => x"204C6F61",
002088 => x"64657220",
002089 => x"77697468",
002090 => x"20444530",
002091 => x"2D4E414E",
002092 => x"4F203332",
002093 => x"4D422073",
002094 => x"7570706F",
002095 => x"72747625",
002096 => x"730A0000",
002097 => x"32303135",
002098 => x"2D31302D",
002099 => x"30330000",
002100 => x"52656164",
002101 => x"790A3E20",
002102 => x"00000000",
002103 => x"3E200000",
002104 => x"454C4600",
002105 => x"4552524F",
002106 => x"523A204E",
002107 => x"6F742061",
002108 => x"6E20454C",
002109 => x"46206669",
002110 => x"6C652E0A",
002111 => x"00000000",
002112 => x"4552524F",
002113 => x"523A2045",
002114 => x"4C462066",
002115 => x"696C6520",
002116 => x"6E6F7420",
002117 => x"74617267",
002118 => x"65747469",
002119 => x"6E672063",
002120 => x"6F727265",
002121 => x"63742070",
002122 => x"726F6365",
002123 => x"73736F72",
002124 => x"20747970",
002125 => x"650A0000",
002126 => x"286E756C",
002127 => x"6C290000",
others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;