-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
--				MEM_SIZE      : natural := 1024;  -- memory cells
--				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				MEM_SIZE      : natural := 2048;  -- memory cells
				LOG2_MEM_SIZE : natural := 11;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
000000 => x"EA000006",
000001 => x"EA0004B5",
000002 => x"EA0004B4",
000003 => x"EA0004B3",
000004 => x"EA0004B2",
000005 => x"EA0004B1",
000006 => x"EA0004B0",
000007 => x"EA0004AF",
000008 => x"E59F0168",
000009 => x"E10F1000",
000010 => x"E3C1107F",
000011 => x"E38110DF",
000012 => x"E129F001",
000013 => x"E1A0D000",
000014 => x"E3A00000",
000015 => x"E1A01000",
000016 => x"E1A02000",
000017 => x"E1A0B000",
000018 => x"E1A07000",
000019 => x"E59FA140",
000020 => x"E1A0E00F",
000021 => x"E1A0F00A",
000022 => x"E3A00003",
000023 => x"E13FF000",
000024 => x"E59FD098",
000025 => x"EB0001EA",
000026 => x"E59F1118",
000027 => x"E59F20B8",
000028 => x"E59F30B8",
000029 => x"E1520003",
000030 => x"0A000002",
000031 => x"E4924004",
000032 => x"E4814004",
000033 => x"EAFFFFFA",
000034 => x"E59F20FC",
000035 => x"E3A03000",
000036 => x"E3A04028",
000037 => x"E4823004",
000038 => x"E2544001",
000039 => x"1AFFFFFC",
000040 => x"E1A04000",
000041 => x"E38443C3",
000042 => x"E3A00000",
000043 => x"E1A0F004",
000044 => x"E92D4000",
000045 => x"E92D1FFF",
000046 => x"E3A04000",
000047 => x"E1A0500D",
000048 => x"E1A0600E",
000049 => x"E59F00CC",
000050 => x"E1A01004",
000051 => x"E4952004",
000052 => x"EB000467",
000053 => x"E354000D",
000054 => x"12844001",
000055 => x"1AFFFFF8",
000056 => x"E59F00B4",
000057 => x"E1A0100D",
000058 => x"EB000461",
000059 => x"E59F00AC",
000060 => x"E2461004",
000061 => x"EB00045E",
000062 => x"E8BD1FFF",
000063 => x"E8FD8000",
000064 => x"007FFFF8",
000065 => x"F0000020",
000066 => x"72253264",
000067 => x"20202530",
000068 => x"38780A00",
000069 => x"73702020",
000070 => x"20253038",
000071 => x"780A0070",
000072 => x"63202020",
000073 => x"25303878",
000074 => x"0A000000",
000075 => x"00010134",
000076 => x"00010184",
000077 => x"00000005",
000078 => x"54410001",
000079 => x"00000001",
000080 => x"00001000",
000081 => x"00000000",
000082 => x"00000004",
000083 => x"54410002",
000084 => x"00800000",
000085 => x"00000000",
000086 => x"00000005",
000087 => x"54410004",
000088 => x"00000001",
000089 => x"000000D0",
000090 => x"00001E00",
000091 => x"00000004",
000092 => x"54410005",
000093 => x"02700000",
000094 => x"00034000",
000095 => x"00000000",
000096 => x"00000000",
000097 => x"00000000",
000098 => x"0007C000",
000099 => x"03F01000",
000100 => x"00002100",
000101 => x"00010814",
000102 => x"00010108",
000103 => x"00010114",
000104 => x"0001011F",
000105 => x"E92D45F0",
000106 => x"E1A04002",
000107 => x"E3A02000",
000108 => x"E5842000",
000109 => x"E1A06001",
000110 => x"E1A0A003",
000111 => x"E0805001",
000112 => x"E1A07002",
000113 => x"E1A08001",
000114 => x"E5D51000",
000115 => x"E59F00CC",
000116 => x"EB000427",
000117 => x"E5D52000",
000118 => x"E2423030",
000119 => x"E3530009",
000120 => x"E2421041",
000121 => x"E3A00000",
000122 => x"8A000006",
000123 => x"E5943000",
000124 => x"E1A03203",
000125 => x"E5843000",
000126 => x"E5D52000",
000127 => x"E0833002",
000128 => x"E2433030",
000129 => x"EA000009",
000130 => x"E3510005",
000131 => x"E2423061",
000132 => x"E3A00000",
000133 => x"8A000007",
000134 => x"E5943000",
000135 => x"E1A03203",
000136 => x"E5843000",
000137 => x"E5D52000",
000138 => x"E0833002",
000139 => x"E2433037",
000140 => x"E5843000",
000141 => x"EA00000B",
000142 => x"E3530005",
000143 => x"E3A00000",
000144 => x"858A7000",
000145 => x"83A00001",
000146 => x"8A000006",
000147 => x"E5943000",
000148 => x"E1A03203",
000149 => x"E5843000",
000150 => x"E5D52000",
000151 => x"E0833002",
000152 => x"E2433057",
000153 => x"EAFFFFF1",
000154 => x"E2883001",
000155 => x"E3570008",
000156 => x"E2855001",
000157 => x"E1A08003",
000158 => x"058A7000",
000159 => x"0A000002",
000160 => x"E3500000",
000161 => x"E2877001",
000162 => x"0AFFFFCE",
000163 => x"E2860001",
000164 => x"E1530000",
000165 => x"D3A00000",
000166 => x"C3A00001",
000167 => x"E8BD85F0",
000168 => x"00011E9C",
000169 => x"E92D4070",
000170 => x"E24DD004",
000171 => x"E1A06002",
000172 => x"E1A0300D",
000173 => x"E1A02001",
000174 => x"E3A01002",
000175 => x"E1A04000",
000176 => x"EBFFFFB7",
000177 => x"E2501000",
000178 => x"E1A0500D",
000179 => x"E1A02006",
000180 => x"E1A00004",
000181 => x"E1A0300D",
000182 => x"0A000003",
000183 => x"E59D1000",
000184 => x"E2811003",
000185 => x"EBFFFFAE",
000186 => x"E1A01000",
000187 => x"E1A00001",
000188 => x"E28DD004",
000189 => x"E8BD8070",
000190 => x"E92D4010",
000191 => x"E1A04000",
000192 => x"EA000000",
000193 => x"EB0003DA",
000194 => x"E2544001",
000195 => x"E59F0004",
000196 => x"2AFFFFFB",
000197 => x"E8BD8010",
000198 => x"00011EA0",
000199 => x"E52DE004",
000200 => x"E59F00CC",
000201 => x"EB0003D2",
000202 => x"E59F00C8",
000203 => x"EB0003D0",
000204 => x"E3A0001D",
000205 => x"EBFFFFEF",
000206 => x"E59F00BC",
000207 => x"EB0003CC",
000208 => x"E59F00B8",
000209 => x"EB0003CA",
000210 => x"E3A00013",
000211 => x"EBFFFFE9",
000212 => x"E59F00AC",
000213 => x"EB0003C6",
000214 => x"E59F00A8",
000215 => x"EB0003C4",
000216 => x"E59F00A4",
000217 => x"EB0003C2",
000218 => x"E3A0001D",
000219 => x"EBFFFFE1",
000220 => x"E59F0098",
000221 => x"EB0003BE",
000222 => x"E59F0094",
000223 => x"EB0003BC",
000224 => x"E3A00013",
000225 => x"EBFFFFDB",
000226 => x"E59F0088",
000227 => x"EB0003B8",
000228 => x"E59F0084",
000229 => x"EB0003B6",
000230 => x"E3A00013",
000231 => x"EBFFFFD5",
000232 => x"E59F0078",
000233 => x"EB0003B2",
000234 => x"E59F0074",
000235 => x"EB0003B0",
000236 => x"E3A00013",
000237 => x"EBFFFFCF",
000238 => x"E59F0068",
000239 => x"EB0003AC",
000240 => x"E59F0064",
000241 => x"EB0003AA",
000242 => x"E3A0001D",
000243 => x"EBFFFFC9",
000244 => x"E59F0058",
000245 => x"EB0003A6",
000246 => x"E59F0054",
000247 => x"EB0003A4",
000248 => x"E3A0000B",
000249 => x"EBFFFFC3",
000250 => x"E59F0048",
000251 => x"E49DE004",
000252 => x"EA00039F",
000253 => x"00011EA4",
000254 => x"00011EB0",
000255 => x"00011EB4",
000256 => x"00011EC8",
000257 => x"00011ED4",
000258 => x"00011EF8",
000259 => x"00011F24",
000260 => x"00011F28",
000261 => x"00011F40",
000262 => x"00011F4C",
000263 => x"00011F78",
000264 => x"00011F84",
000265 => x"00011FA8",
000266 => x"00011FB4",
000267 => x"00011FC0",
000268 => x"00011FC4",
000269 => x"00011FD4",
000270 => x"00011FE8",
000271 => x"E92D4010",
000272 => x"E1A01000",
000273 => x"E1A04000",
000274 => x"E59F0014",
000275 => x"EB000388",
000276 => x"E59F0010",
000277 => x"E5942000",
000278 => x"E1A01004",
000279 => x"E8BD4010",
000280 => x"EA000383",
000281 => x"00011FF8",
000282 => x"00012008",
000283 => x"E2400001",
000284 => x"E92D4010",
000285 => x"E1A04001",
000286 => x"E3500004",
000287 => x"979FF100",
000288 => x"EA000039",
000289 => x"00010498",
000290 => x"000104D8",
000291 => x"000104EC",
000292 => x"00010518",
000293 => x"0001053C",
000294 => x"E59F10EC",
000295 => x"E59F00EC",
000296 => x"EB000373",
000297 => x"E3A01602",
000298 => x"E3A00505",
000299 => x"EB00015B",
000300 => x"E3500602",
000301 => x"E1A04000",
000302 => x"81A01000",
000303 => x"8A000027",
000304 => x"E59F00CC",
000305 => x"EB00036A",
000306 => x"E1A01004",
000307 => x"E3A00505",
000308 => x"E8BD4010",
000309 => x"EA0001F7",
000310 => x"EBFFFF8F",
000311 => x"EBFFFEF3",
000312 => x"E3A00010",
000313 => x"EBFFFF83",
000314 => x"EA000008",
000315 => x"E3A01702",
000316 => x"E59F00A0",
000317 => x"EB00035E",
000318 => x"E3A00010",
000319 => x"EBFFFF7D",
000320 => x"E59F0094",
000321 => x"EB00035A",
000322 => x"E3A00702",
000323 => x"EBFFFED5",
000324 => x"E8BD4010",
000325 => x"EA000374",
000326 => x"E3A01901",
000327 => x"E59F0074",
000328 => x"EB000353",
000329 => x"E3A00010",
000330 => x"EBFFFF72",
000331 => x"E59F0068",
000332 => x"EB00034F",
000333 => x"E3A00901",
000334 => x"EAFFFFF3",
000335 => x"E59F1048",
000336 => x"E59F0048",
000337 => x"EB00034A",
000338 => x"E1A00004",
000339 => x"E3A01602",
000340 => x"EB000132",
000341 => x"E3500602",
000342 => x"98BD8010",
000343 => x"E1A01000",
000344 => x"E59F0038",
000345 => x"E8BD4010",
000346 => x"EA000341",
000347 => x"E59F0024",
000348 => x"EB00033F",
000349 => x"E3A00010",
000350 => x"EBFFFF5E",
000351 => x"E59F0018",
000352 => x"EB00033B",
000353 => x"E1A00004",
000354 => x"EAFFFFDF",
000355 => x"00012024",
000356 => x"00012020",
000357 => x"00012084",
000358 => x"00012090",
000359 => x"00012004",
000360 => x"00012064",
000361 => x"E92D4010",
000362 => x"E59F3250",
000363 => x"E5D0C001",
000364 => x"E1A0E000",
000365 => x"E893000F",
000366 => x"E24DD020",
000367 => x"E35C0000",
000368 => x"E1A0400D",
000369 => x"E88D000F",
000370 => x"0A00008A",
000371 => x"E35C000D",
000372 => x"1A000011",
000373 => x"E5DE0000",
000374 => x"E350006C",
000375 => x"0A000005",
000376 => x"E3500073",
000377 => x"0A000006",
000378 => x"E3500068",
000379 => x"1A00000C",
000380 => x"EBFFFF49",
000381 => x"EA00007F",
000382 => x"E3A00001",
000383 => x"E3A01000",
000384 => x"EA000034",
000385 => x"EBFFFEA9",
000386 => x"E3A00010",
000387 => x"EBFFFF39",
000388 => x"E59F01EC",
000389 => x"EB000316",
000390 => x"EA000076",
000391 => x"E35C0020",
000392 => x"0A000002",
000393 => x"E59F01DC",
000394 => x"E1A0100D",
000395 => x"EA000070",
000396 => x"E5DE3000",
000397 => x"E353006A",
000398 => x"0A00001D",
000399 => x"8A000004",
000400 => x"E3530062",
000401 => x"0A00004D",
000402 => x"E3530064",
000403 => x"1A000066",
000404 => x"EA000006",
000405 => x"E3530072",
000406 => x"0A000040",
000407 => x"E3530077",
000408 => x"0A00004F",
000409 => x"E3530070",
000410 => x"1A00005F",
000411 => x"EA00001B",
000412 => x"E1A0000E",
000413 => x"E28D1010",
000414 => x"E28D2014",
000415 => x"EBFFFF08",
000416 => x"E3500000",
000417 => x"159D4010",
000418 => x"1A000001",
000419 => x"EA000059",
000420 => x"EBFFFF69",
000421 => x"E59D3010",
000422 => x"E59D2014",
000423 => x"E0833002",
000424 => x"E1540003",
000425 => x"E1A00004",
000426 => x"E2844004",
000427 => x"3AFFFFF7",
000428 => x"EA000050",
000429 => x"E1A0000E",
000430 => x"E3A01002",
000431 => x"E28D2010",
000432 => x"E28D3018",
000433 => x"EBFFFEB6",
000434 => x"E3500000",
000435 => x"0A000049",
000436 => x"E3A00000",
000437 => x"E59D1010",
000438 => x"EBFFFF63",
000439 => x"EA000045",
000440 => x"E1A0000E",
000441 => x"E3A01002",
000442 => x"E28D2010",
000443 => x"E28D3018",
000444 => x"EBFFFEAB",
000445 => x"E3500000",
000446 => x"0A00003E",
000447 => x"E3A03000",
000448 => x"E58D3018",
000449 => x"E59D3010",
000450 => x"E4D34001",
000451 => x"E58D3010",
000452 => x"EA00000B",
000453 => x"E3540000",
000454 => x"0A000003",
000455 => x"EB0002F6",
000456 => x"E354000D",
000457 => x"E59F00D8",
000458 => x"0B0002D1",
000459 => x"E59D2010",
000460 => x"E59D3018",
000461 => x"E4D24001",
000462 => x"E2833001",
000463 => x"E58D2010",
000464 => x"E58D3018",
000465 => x"E3140080",
000466 => x"E1A00004",
000467 => x"1A000029",
000468 => x"E59D3018",
000469 => x"E3530A01",
000470 => x"3AFFFFED",
000471 => x"EA000025",
000472 => x"E1A0000E",
000473 => x"E3A01002",
000474 => x"E28D2010",
000475 => x"E28D3018",
000476 => x"EBFFFE8B",
000477 => x"E3500000",
000478 => x"0A00001E",
000479 => x"EA000017",
000480 => x"E1A0000E",
000481 => x"E3A01002",
000482 => x"E28D2010",
000483 => x"E28D3018",
000484 => x"EBFFFE83",
000485 => x"E3500000",
000486 => x"13A00005",
000487 => x"1AFFFFCC",
000488 => x"EA000014",
000489 => x"E1A0000E",
000490 => x"E28D1010",
000491 => x"E28D201C",
000492 => x"EBFFFEBB",
000493 => x"E3500000",
000494 => x"0A00000E",
000495 => x"E59D1010",
000496 => x"E59F0044",
000497 => x"EB0002AA",
000498 => x"E59D101C",
000499 => x"E59F003C",
000500 => x"EB0002A7",
000501 => x"E59D201C",
000502 => x"E59D3010",
000503 => x"E5832000",
000504 => x"E59D0010",
000505 => x"EBFFFF14",
000506 => x"EA000002",
000507 => x"E59F0014",
000508 => x"E1A0100D",
000509 => x"EB00029E",
000510 => x"E28DD020",
000511 => x"E8BD8010",
000512 => x"000120A8",
000513 => x"00012004",
000514 => x"00012020",
000515 => x"00011FF8",
000516 => x"0001209C",
000517 => x"E92D41F0",
000518 => x"E3A0100C",
000519 => x"E24DD028",
000520 => x"E59F2170",
000521 => x"E59F0170",
000522 => x"EB000291",
000523 => x"EBFFFEBA",
000524 => x"E59F0168",
000525 => x"EB00028E",
000526 => x"E3A06000",
000527 => x"E1A07006",
000528 => x"E1A08006",
000529 => x"EA000001",
000530 => x"E1A06008",
000531 => x"E3A07000",
000532 => x"E3A00FFA",
000533 => x"EB0002B0",
000534 => x"E2504000",
000535 => x"BAFFFFFB",
000536 => x"E354001B",
000537 => x"0A00001C",
000538 => x"E3570001",
000539 => x"0354005B",
000540 => x"13A05000",
000541 => x"03A05001",
000542 => x"03A07002",
000543 => x"0A00001D",
000544 => x"E3570002",
000545 => x"1A000038",
000546 => x"E3540041",
000547 => x"01A04005",
000548 => x"11A07005",
000549 => x"1AFFFFED",
000550 => x"EA000000",
000551 => x"EB000296",
000552 => x"E1540006",
000553 => x"E3A00008",
000554 => x"E2844001",
000555 => x"BAFFFFFA",
000556 => x"E3A04000",
000557 => x"EA000005",
000558 => x"E28D3014",
000559 => x"E7D42003",
000560 => x"E1A00002",
000561 => x"E7C4200D",
000562 => x"EB00028B",
000563 => x"E2844001",
000564 => x"E1540008",
000565 => x"BAFFFFF7",
000566 => x"EAFFFFDA",
000567 => x"E3A07001",
000568 => x"EA000004",
000569 => x"E28D2028",
000570 => x"E0823006",
000571 => x"E5434028",
000572 => x"E2866001",
000573 => x"E3A07000",
000574 => x"E3560012",
000575 => x"D3A03000",
000576 => x"C3A03001",
000577 => x"E354000D",
000578 => x"03833001",
000579 => x"E3530000",
000580 => x"0AFFFFCE",
000581 => x"E3560001",
000582 => x"DA000007",
000583 => x"E3A01000",
000584 => x"E7D1200D",
000585 => x"E28D3014",
000586 => x"E7C12003",
000587 => x"E2811001",
000588 => x"E3510014",
000589 => x"1AFFFFF9",
000590 => x"E2468001",
000591 => x"E28D2028",
000592 => x"E0823006",
000593 => x"E3A04000",
000594 => x"E5434028",
000595 => x"E59F0050",
000596 => x"EB000247",
000597 => x"E1A0000D",
000598 => x"EBFFFF11",
000599 => x"E59F0044",
000600 => x"EB000243",
000601 => x"E1A06004",
000602 => x"EAFFFFB8",
000603 => x"EB000262",
000604 => x"E3540008",
000605 => x"13A03000",
000606 => x"03A03001",
000607 => x"E3560000",
000608 => x"D3A03000",
000609 => x"E3530000",
000610 => x"12466001",
000611 => x"11A07005",
000612 => x"1AFFFFD8",
000613 => x"EAFFFFD2",
000614 => x"000120EC",
000615 => x"000120B8",
000616 => x"000120F8",
000617 => x"00012004",
000618 => x"00012104",
000619 => x"E92D4010",
000620 => x"E3A0C000",
000621 => x"E1A04000",
000622 => x"E1A0E00C",
000623 => x"E1A00001",
000624 => x"EA00000A",
000625 => x"E7DE3004",
000626 => x"E023342C",
000627 => x"E1A03083",
000628 => x"E0832001",
000629 => x"E7D31001",
000630 => x"E5D23001",
000631 => x"E1833401",
000632 => x"E023340C",
000633 => x"E1A03803",
000634 => x"E28EE001",
000635 => x"E1A0C823",
000636 => x"E15E0000",
000637 => x"E59F1008",
000638 => x"BAFFFFF1",
000639 => x"E1A0000C",
000640 => x"E8BD8010",
000641 => x"00011C9C",
000642 => x"E52DE004",
000643 => x"E3A00F4B",
000644 => x"EB000241",
000645 => x"E3500000",
000646 => x"AAFFFFFB",
000647 => x"E49DF004",
000648 => x"E92D4FF0",
000649 => x"E3A07000",
000650 => x"E24DDB01",
000651 => x"E24DD008",
000652 => x"E1A0B000",
000653 => x"E1A09001",
000654 => x"E3A0A019",
000655 => x"E3A04043",
000656 => x"E3A08001",
000657 => x"E1A06007",
000658 => x"EA000000",
000659 => x"E3A04015",
000660 => x"E3A05000",
000661 => x"E3540000",
000662 => x"11A00004",
000663 => x"1B000226",
000664 => x"E3A00FFA",
000665 => x"EB00022C",
000666 => x"E3500000",
000667 => x"BA000019",
000668 => x"E3500002",
000669 => x"0A000025",
000670 => x"CA000002",
000671 => x"E3500001",
000672 => x"1A000014",
000673 => x"EA000004",
000674 => x"E3500004",
000675 => x"0A000004",
000676 => x"E3500018",
000677 => x"1A00000F",
000678 => x"EA000005",
000679 => x"E3A05080",
000680 => x"EA00001B",
000681 => x"E3A00006",
000682 => x"EB000213",
000683 => x"EBFFFFD5",
000684 => x"EA00007C",
000685 => x"E3A00FFA",
000686 => x"EB000217",
000687 => x"E3500018",
000688 => x"1A000004",
000689 => x"EBFFFFCF",
000690 => x"E3A00006",
000691 => x"EB00020A",
000692 => x"E3E06000",
000693 => x"EA000073",
000694 => x"E2855001",
000695 => x"E3550050",
000696 => x"1AFFFFDB",
000697 => x"E3540043",
000698 => x"0AFFFFD7",
000699 => x"EBFFFFC5",
000700 => x"E3A00018",
000701 => x"EB000200",
000702 => x"E3A00018",
000703 => x"EB0001FE",
000704 => x"E3A00018",
000705 => x"EB0001FC",
000706 => x"E3E06001",
000707 => x"EA000065",
000708 => x"E3A05B01",
000709 => x"E3540043",
000710 => x"03A07001",
000711 => x"E1A00000",
000712 => x"E5CD0002",
000713 => x"E1A00000",
000714 => x"E3A04000",
000715 => x"EA000006",
000716 => x"EB0001F9",
000717 => x"E28D3008",
000718 => x"E3500000",
000719 => x"E2433006",
000720 => x"E2844001",
000721 => x"BA000052",
000722 => x"E7C40003",
000723 => x"E3570000",
000724 => x"13A03004",
000725 => x"03A03003",
000726 => x"E0853003",
000727 => x"E1540003",
000728 => x"E3A00FFA",
000729 => x"BAFFFFF1",
000730 => x"E5DD3004",
000731 => x"E5DD2003",
000732 => x"E1E03003",
000733 => x"E20330FF",
000734 => x"E1520003",
000735 => x"1A000044",
000736 => x"E1520008",
000737 => x"0A000002",
000738 => x"E2483001",
000739 => x"E1520003",
000740 => x"1A00003F",
000741 => x"E3570000",
000742 => x"E28D4008",
000743 => x"E2444006",
000744 => x"01A01007",
000745 => x"02840003",
000746 => x"01A02001",
000747 => x"0A00000D",
000748 => x"E2840003",
000749 => x"E1A01005",
000750 => x"EBFFFF7B",
000751 => x"E0843005",
000752 => x"E5D32004",
000753 => x"E5D33003",
000754 => x"E0822403",
000755 => x"E1A02802",
000756 => x"E1500822",
000757 => x"1A00002E",
000758 => x"EA00000C",
000759 => x"E5503001",
000760 => x"E0813003",
000761 => x"E20310FF",
000762 => x"E1520005",
000763 => x"E2800001",
000764 => x"E2822001",
000765 => x"BAFFFFF8",
000766 => x"E28D2B01",
000767 => x"E2822008",
000768 => x"E0823005",
000769 => x"E5533403",
000770 => x"E1530001",
000771 => x"1A000020",
000772 => x"E5DD3003",
000773 => x"E1530008",
000774 => x"1A00000F",
000775 => x"E0663009",
000776 => x"E1550003",
000777 => x"B1A04005",
000778 => x"A1A04003",
000779 => x"E3540000",
000780 => x"DA000005",
000781 => x"E28D1008",
000782 => x"E08B0006",
000783 => x"E2411003",
000784 => x"E1A02004",
000785 => x"EB0002C5",
000786 => x"E0866004",
000787 => x"E2883001",
000788 => x"E20380FF",
000789 => x"E3A0A019",
000790 => x"EA00000B",
000791 => x"E24AA001",
000792 => x"E35A0000",
000793 => x"CA000008",
000794 => x"EBFFFF66",
000795 => x"E3A00018",
000796 => x"EB0001A1",
000797 => x"E3A00018",
000798 => x"EB00019F",
000799 => x"E3A00018",
000800 => x"EB00019D",
000801 => x"E3E06002",
000802 => x"EA000006",
000803 => x"E3A00006",
000804 => x"EA000001",
000805 => x"EBFFFF5B",
000806 => x"E3A00015",
000807 => x"EB000196",
000808 => x"E3A04000",
000809 => x"EAFFFF69",
000810 => x"E1A00006",
000811 => x"E28DD008",
000812 => x"E28DDB01",
000813 => x"E8BD8FF0",
000814 => x"E92D40F0",
000815 => x"E1A05000",
000816 => x"E2804012",
000817 => x"E59F01BC",
000818 => x"EB000169",
000819 => x"E5D53012",
000820 => x"E5D41001",
000821 => x"E59F01B0",
000822 => x"E1811403",
000823 => x"EB000164",
000824 => x"E2850001",
000825 => x"E59F11A4",
000826 => x"E3A02003",
000827 => x"EB000287",
000828 => x"E2506000",
000829 => x"159F0198",
000830 => x"1A000005",
000831 => x"E5D43001",
000832 => x"E5D52012",
000833 => x"E1833402",
000834 => x"E3530028",
000835 => x"0A000003",
000836 => x"E59F0180",
000837 => x"EB000156",
000838 => x"E3A00001",
000839 => x"E8BD80F0",
000840 => x"E5D5302C",
000841 => x"E5D5102D",
000842 => x"E59F016C",
000843 => x"E1811403",
000844 => x"EB00014F",
000845 => x"E1A04006",
000846 => x"EA00000A",
000847 => x"E5D5102A",
000848 => x"E595201C",
000849 => x"E5D5302B",
000850 => x"E0852002",
000851 => x"E1833401",
000852 => x"E0232394",
000853 => x"E5932014",
000854 => x"E5931008",
000855 => x"E0811002",
000856 => x"EB000143",
000857 => x"E2844001",
000858 => x"E5D5202C",
000859 => x"E5D5302D",
000860 => x"E1833402",
000861 => x"E1540003",
000862 => x"E59F0120",
000863 => x"3AFFFFEE",
000864 => x"E3A07000",
000865 => x"EA000038",
000866 => x"E5952020",
000867 => x"E5D5102E",
000868 => x"E5D5302F",
000869 => x"E0852002",
000870 => x"E1833401",
000871 => x"E0242397",
000872 => x"E5943004",
000873 => x"E3530001",
000874 => x"1A000018",
000875 => x"E5943014",
000876 => x"E3530000",
000877 => x"0A00002B",
000878 => x"E594300C",
000879 => x"E3530000",
000880 => x"13A06000",
000881 => x"1A00000E",
000882 => x"EA000026",
000883 => x"E5942010",
000884 => x"E0862002",
000885 => x"E0851002",
000886 => x"E5D13002",
000887 => x"E5D10003",
000888 => x"E7D5C002",
000889 => x"E1A03803",
000890 => x"E5D12001",
000891 => x"E1833C00",
000892 => x"E594E00C",
000893 => x"E183300C",
000894 => x"E1833402",
000895 => x"E78E3006",
000896 => x"E2866004",
000897 => x"E5943014",
000898 => x"E1560003",
000899 => x"3AFFFFEE",
000900 => x"E5943004",
000901 => x"E3530008",
000902 => x"1A000012",
000903 => x"E5943014",
000904 => x"E3530000",
000905 => x"0A00000F",
000906 => x"E594300C",
000907 => x"E3530000",
000908 => x"15941010",
000909 => x"1A000006",
000910 => x"EA00000A",
000911 => x"E594300C",
000912 => x"E0813003",
000913 => x"E0623003",
000914 => x"E3A02000",
000915 => x"E5832000",
000916 => x"E2811004",
000917 => x"E2842010",
000918 => x"E892000C",
000919 => x"E0823003",
000920 => x"E1510003",
000921 => x"3AFFFFF4",
000922 => x"E2877001",
000923 => x"E5D52030",
000924 => x"E5D53031",
000925 => x"E1833402",
000926 => x"E1570003",
000927 => x"3AFFFFC1",
000928 => x"E3A00000",
000929 => x"E8BD80F0",
000930 => x"00012108",
000931 => x"0001211C",
000932 => x"00012140",
000933 => x"00012144",
000934 => x"00012160",
000935 => x"00012198",
000936 => x"000121B8",
000937 => x"E5903000",
000938 => x"E20110FF",
000939 => x"E3530000",
000940 => x"14C31001",
000941 => x"E1A02000",
000942 => x"E1A00001",
000943 => x"15823000",
000944 => x"11A0F00E",
000945 => x"EA00010C",
000946 => x"E92D45F0",
000947 => x"E2525000",
000948 => x"E1A08000",
000949 => x"E1A07001",
000950 => x"C3A02000",
000951 => x"CA000001",
000952 => x"EA000009",
000953 => x"E2822001",
000954 => x"E7D21007",
000955 => x"E3510000",
000956 => x"1AFFFFFB",
000957 => x"E1520005",
000958 => x"A1A05001",
000959 => x"B0625005",
000960 => x"E3130002",
000961 => x"13A0A030",
000962 => x"1A000000",
000963 => x"E3A0A020",
000964 => x"E3130001",
000965 => x"13A06000",
000966 => x"01A04005",
000967 => x"0A000002",
000968 => x"EA00000A",
000969 => x"EBFFFFDE",
000970 => x"E2444001",
000971 => x"E3540000",
000972 => x"E1A00008",
000973 => x"E20A10FF",
000974 => x"CAFFFFF9",
000975 => x"E0646005",
000976 => x"E1A05004",
000977 => x"EA000001",
000978 => x"EBFFFFD5",
000979 => x"E2866001",
000980 => x"E5D73000",
000981 => x"E2531000",
000982 => x"E1A00008",
000983 => x"E2877001",
000984 => x"1AFFFFF8",
000985 => x"EA000001",
000986 => x"EBFFFFCD",
000987 => x"E2866001",
000988 => x"E3550000",
000989 => x"E1A00008",
000990 => x"E20A10FF",
000991 => x"E2455001",
000992 => x"CAFFFFF8",
000993 => x"E1A00006",
000994 => x"E8BD85F0",
000995 => x"E92D4FF0",
000996 => x"E2514000",
000997 => x"E24DD010",
000998 => x"E1A05002",
000999 => x"E1A09000",
001000 => x"E28D6034",
001001 => x"E8960C40",
001002 => x"1A000007",
001003 => x"E3A0C030",
001004 => x"E1A02006",
001005 => x"E1A0300A",
001006 => x"E1A0100D",
001007 => x"E5CDC000",
001008 => x"E5CD4001",
001009 => x"EBFFFFBF",
001010 => x"EA00003C",
001011 => x"E2533000",
001012 => x"13A03001",
001013 => x"E352000A",
001014 => x"13A03000",
001015 => x"E3530000",
001016 => x"0A000003",
001017 => x"E3540000",
001018 => x"B2644000",
001019 => x"B3A08001",
001020 => x"BA000000",
001021 => x"E3A08000",
001022 => x"E3A03000",
001023 => x"E28D700F",
001024 => x"E5CD300F",
001025 => x"EA000010",
001026 => x"E3550010",
001027 => x"0A000002",
001028 => x"EB0000CD",
001029 => x"E0030095",
001030 => x"E0633004",
001031 => x"E3530009",
001032 => x"E083200B",
001033 => x"C242303A",
001034 => x"E2833030",
001035 => x"E3550010",
001036 => x"E1A00004",
001037 => x"E1A01005",
001038 => x"E5673001",
001039 => x"01A04224",
001040 => x"0A000001",
001041 => x"EB0000C0",
001042 => x"E1A04000",
001043 => x"E3540000",
001044 => x"E1A00004",
001045 => x"E1A01005",
001046 => x"E204300F",
001047 => x"1AFFFFE9",
001048 => x"E3580000",
001049 => x"E1A02007",
001050 => x"01A04008",
001051 => x"0A00000D",
001052 => x"E3560000",
001053 => x"0A000007",
001054 => x"E31A0002",
001055 => x"0A000005",
001056 => x"E1A00009",
001057 => x"E3A0102D",
001058 => x"EBFFFF85",
001059 => x"E2466001",
001060 => x"E3A04001",
001061 => x"EA000003",
001062 => x"E3A0302D",
001063 => x"E5423001",
001064 => x"E2477001",
001065 => x"E3A04000",
001066 => x"E1A00009",
001067 => x"E1A01007",
001068 => x"E1A02006",
001069 => x"E1A0300A",
001070 => x"EBFFFF82",
001071 => x"E0840000",
001072 => x"E28DD010",
001073 => x"E8BD8FF0",
001074 => x"E92D41F0",
001075 => x"E1A07000",
001076 => x"E24DD010",
001077 => x"E1A04001",
001078 => x"E1A05002",
001079 => x"E3A06000",
001080 => x"EA00005C",
001081 => x"E3530025",
001082 => x"1A000051",
001083 => x"E5F43001",
001084 => x"E3530000",
001085 => x"0A00005A",
001086 => x"E3530025",
001087 => x"0A000050",
001088 => x"E353002D",
001089 => x"13A08000",
001090 => x"02844001",
001091 => x"03A08001",
001092 => x"EA000001",
001093 => x"E2844001",
001094 => x"E3888002",
001095 => x"E5D43000",
001096 => x"E3530030",
001097 => x"0AFFFFFA",
001098 => x"E3A0E000",
001099 => x"EA000003",
001100 => x"E3A0300A",
001101 => x"E023239E",
001102 => x"E2844001",
001103 => x"E243E030",
001104 => x"E5D42000",
001105 => x"E2423030",
001106 => x"E3530009",
001107 => x"9AFFFFF7",
001108 => x"E3520073",
001109 => x"1A000007",
001110 => x"E4953004",
001111 => x"E59F110C",
001112 => x"E3530000",
001113 => x"11A01003",
001114 => x"E1A0200E",
001115 => x"E1A03008",
001116 => x"E1A00007",
001117 => x"EA00002C",
001118 => x"E3520064",
001119 => x"1A00000A",
001120 => x"E4951004",
001121 => x"E1A00007",
001122 => x"E3A0200A",
001123 => x"E3A03001",
001124 => x"E58DE000",
001125 => x"E58D8004",
001126 => x"E3A0C061",
001127 => x"E58DC008",
001128 => x"EBFFFF79",
001129 => x"E0866000",
001130 => x"EA000029",
001131 => x"E3520078",
001132 => x"04951004",
001133 => x"01A00007",
001134 => x"03A02010",
001135 => x"0A00000E",
001136 => x"E3520058",
001137 => x"1A000007",
001138 => x"E4951004",
001139 => x"E1A00007",
001140 => x"E3A02010",
001141 => x"E3A03000",
001142 => x"E3A0C041",
001143 => x"E58DE000",
001144 => x"E58D8004",
001145 => x"EAFFFFEC",
001146 => x"E3520075",
001147 => x"1A000004",
001148 => x"E4951004",
001149 => x"E1A00007",
001150 => x"E3A0200A",
001151 => x"E3A03000",
001152 => x"EAFFFFE2",
001153 => x"E3520063",
001154 => x"1A000011",
001155 => x"E495C004",
001156 => x"E5CDC00E",
001157 => x"E3A0C000",
001158 => x"E5CDC00F",
001159 => x"E1A0200E",
001160 => x"E1A03008",
001161 => x"E1A00007",
001162 => x"E28D100E",
001163 => x"EBFFFF25",
001164 => x"EAFFFFDB",
001165 => x"E353000A",
001166 => x"01A00007",
001167 => x"03A0100D",
001168 => x"0BFFFF17",
001169 => x"E1A00007",
001170 => x"E5D41000",
001171 => x"EBFFFF14",
001172 => x"E2866001",
001173 => x"E2844001",
001174 => x"E5D43000",
001175 => x"E3530000",
001176 => x"1AFFFF9F",
001177 => x"E1A00006",
001178 => x"E28DD010",
001179 => x"E8BD81F0",
001180 => x"000121D4",
001181 => x"E92D000F",
001182 => x"E52DE004",
001183 => x"E24DD004",
001184 => x"E28D0004",
001185 => x"E3A03000",
001186 => x"E5203004",
001187 => x"E59D1008",
001188 => x"E1A0000D",
001189 => x"E28D200C",
001190 => x"EBFFFF8A",
001191 => x"E28DD004",
001192 => x"E49DE004",
001193 => x"E28DD010",
001194 => x"E1A0F00E",
001195 => x"E92D000E",
001196 => x"E52DE004",
001197 => x"E24DD004",
001198 => x"E28D3004",
001199 => x"E5230004",
001200 => x"E59D1008",
001201 => x"E1A0000D",
001202 => x"E28D200C",
001203 => x"EBFFFF7D",
001204 => x"E28DD004",
001205 => x"E49DE004",
001206 => x"E28DD00C",
001207 => x"E1A0F00E",
001208 => x"E59FB46C",
001209 => x"E58B0000",
001210 => x"EAFFFFFC",
001211 => x"E59FB460",
001212 => x"E3A0A011",
001213 => x"E58BA000",
001214 => x"EAFFFFFB",
001215 => x"E59F1454",
001216 => x"E59F3454",
001217 => x"E5932000",
001218 => x"E2022020",
001219 => x"E3520000",
001220 => x"05810000",
001221 => x"01B0F00E",
001222 => x"1AFFFFF9",
001223 => x"E59F2434",
001224 => x"E59F3434",
001225 => x"E1A01580",
001226 => x"E0811480",
001227 => x"E5930000",
001228 => x"E2100010",
001229 => x"05920000",
001230 => x"01A0F00E",
001231 => x"E2511001",
001232 => x"1AFFFFF9",
001233 => x"E3E00000",
001234 => x"E1B0F00E",
001235 => x"E92D4010",
001236 => x"E2002102",
001237 => x"E2013102",
001238 => x"E0224003",
001239 => x"E3100102",
001240 => x"11E00000",
001241 => x"12800001",
001242 => x"E3110102",
001243 => x"11E01001",
001244 => x"12811001",
001245 => x"E1A02001",
001246 => x"E1A01000",
001247 => x"E3520000",
001248 => x"0A000011",
001249 => x"E3A00000",
001250 => x"E3A03001",
001251 => x"E3530000",
001252 => x"03A03201",
001253 => x"0A000003",
001254 => x"E1520001",
001255 => x"91A02082",
001256 => x"91A03083",
001257 => x"9AFFFFF8",
001258 => x"E1510002",
001259 => x"20411002",
001260 => x"20800003",
001261 => x"E1B030A3",
001262 => x"31A020A2",
001263 => x"3AFFFFF9",
001264 => x"E3140102",
001265 => x"11E00000",
001266 => x"12800001",
001267 => x"E8FD8010",
001268 => x"E92D4070",
001269 => x"E1A06000",
001270 => x"E1862001",
001271 => x"E3120003",
001272 => x"1A00002A",
001273 => x"E8B1003C",
001274 => x"E31200FF",
001275 => x"13120CFF",
001276 => x"131208FF",
001277 => x"131204FF",
001278 => x"14862004",
001279 => x"02411004",
001280 => x"131300FF",
001281 => x"13130CFF",
001282 => x"131308FF",
001283 => x"131304FF",
001284 => x"14863004",
001285 => x"02411004",
001286 => x"131400FF",
001287 => x"13140CFF",
001288 => x"131408FF",
001289 => x"131404FF",
001290 => x"14864004",
001291 => x"02411004",
001292 => x"131500FF",
001293 => x"13150CFF",
001294 => x"131508FF",
001295 => x"131504FF",
001296 => x"14865004",
001297 => x"02411004",
001298 => x"1AFFFFE5",
001299 => x"E4913004",
001300 => x"E4C63001",
001301 => x"E21340FF",
001302 => x"08FD8070",
001303 => x"E1A03423",
001304 => x"E4C63001",
001305 => x"E21340FF",
001306 => x"08FD8070",
001307 => x"E1A03423",
001308 => x"E4C63001",
001309 => x"E21340FF",
001310 => x"08FD8070",
001311 => x"E1A03423",
001312 => x"E4C63001",
001313 => x"E21340FF",
001314 => x"08FD8070",
001315 => x"EAFFFFEE",
001316 => x"E4D13001",
001317 => x"E4C63001",
001318 => x"E3530000",
001319 => x"08FD8070",
001320 => x"E4D13001",
001321 => x"E4C63001",
001322 => x"E3530000",
001323 => x"08FD8070",
001324 => x"E4D13001",
001325 => x"E4C63001",
001326 => x"E3530000",
001327 => x"08FD8070",
001328 => x"E4D13001",
001329 => x"E4C63001",
001330 => x"E3530000",
001331 => x"08FD8070",
001332 => x"EAFFFFEE",
001333 => x"E92D41F0",
001334 => x"E1802001",
001335 => x"E3120003",
001336 => x"1A000018",
001337 => x"E8B0001C",
001338 => x"E8B100E0",
001339 => x"E1520005",
001340 => x"1A000012",
001341 => x"01530006",
001342 => x"1A00002B",
001343 => x"01540007",
001344 => x"1A000049",
001345 => x"E31200FF",
001346 => x"13120CFF",
001347 => x"131208FF",
001348 => x"131204FF",
001349 => x"131300FF",
001350 => x"13130CFF",
001351 => x"131308FF",
001352 => x"131304FF",
001353 => x"131400FF",
001354 => x"13140CFF",
001355 => x"131408FF",
001356 => x"131404FF",
001357 => x"1AFFFFEA",
001358 => x"03A00000",
001359 => x"08FD81F0",
001360 => x"E240000C",
001361 => x"E241100C",
001362 => x"E4D02001",
001363 => x"E4D13001",
001364 => x"E0324003",
001365 => x"1A00005A",
001366 => x"E4D05001",
001367 => x"E4D16001",
001368 => x"E3520000",
001369 => x"0A000054",
001370 => x"E0357006",
001371 => x"1A000054",
001372 => x"E4D02001",
001373 => x"E4D13001",
001374 => x"E3550000",
001375 => x"0A00004E",
001376 => x"E0324003",
001377 => x"1A00004E",
001378 => x"E4D05001",
001379 => x"E4D16001",
001380 => x"E3520000",
001381 => x"0A000048",
001382 => x"E0357006",
001383 => x"1A000048",
001384 => x"E3550000",
001385 => x"0A000044",
001386 => x"1AFFFFE6",
001387 => x"E31200FF",
001388 => x"13120CFF",
001389 => x"131208FF",
001390 => x"131204FF",
001391 => x"0A00003E",
001392 => x"E2400008",
001393 => x"E2411008",
001394 => x"E4D02001",
001395 => x"E4D13001",
001396 => x"E0324003",
001397 => x"1A00003A",
001398 => x"E4D05001",
001399 => x"E4D16001",
001400 => x"E3520000",
001401 => x"0A000034",
001402 => x"E0357006",
001403 => x"1A000034",
001404 => x"E4D02001",
001405 => x"E4D13001",
001406 => x"E3550000",
001407 => x"0A00002E",
001408 => x"E0324003",
001409 => x"1A00002E",
001410 => x"E4D05001",
001411 => x"E4D16001",
001412 => x"E3520000",
001413 => x"0A000028",
001414 => x"E0357006",
001415 => x"1A000028",
001416 => x"E3550000",
001417 => x"0A000024",
001418 => x"1AFFFFC6",
001419 => x"E31200FF",
001420 => x"13120CFF",
001421 => x"131208FF",
001422 => x"131204FF",
001423 => x"131300FF",
001424 => x"13130CFF",
001425 => x"131308FF",
001426 => x"131304FF",
001427 => x"0A00001A",
001428 => x"E2400004",
001429 => x"E2411004",
001430 => x"E4D02001",
001431 => x"E4D13001",
001432 => x"E0324003",
001433 => x"1A000016",
001434 => x"E4D05001",
001435 => x"E4D16001",
001436 => x"E3520000",
001437 => x"0A000010",
001438 => x"E0357006",
001439 => x"1A000010",
001440 => x"E4D02001",
001441 => x"E4D13001",
001442 => x"E3550000",
001443 => x"0A00000A",
001444 => x"E0324003",
001445 => x"1A00000A",
001446 => x"E4D05001",
001447 => x"E4D16001",
001448 => x"E3520000",
001449 => x"0A000004",
001450 => x"E0357006",
001451 => x"1A000004",
001452 => x"E3550000",
001453 => x"0A000000",
001454 => x"1AFFFFA2",
001455 => x"03A00000",
001456 => x"08FD81F0",
001457 => x"E0450006",
001458 => x"E8FD81F0",
001459 => x"E59F107C",
001460 => x"E5811000",
001461 => x"E1A0F00E",
001462 => x"E59F1070",
001463 => x"E5910000",
001464 => x"E2800801",
001465 => x"E5810000",
001466 => x"E1A0F00E",
001467 => x"E92D4010",
001468 => x"E3520000",
001469 => x"0A000004",
001470 => x"E0804002",
001471 => x"E4D13001",
001472 => x"E4C03001",
001473 => x"E1500004",
001474 => x"1AFFFFFB",
001475 => x"E8FD8010",
001476 => x"E92D4070",
001477 => x"E3520000",
001478 => x"03A00001",
001479 => x"0A00000A",
001480 => x"E3A03000",
001481 => x"E2833001",
001482 => x"E4D04001",
001483 => x"E4D15001",
001484 => x"E0546005",
001485 => x"11A00006",
001486 => x"1A000003",
001487 => x"E1530002",
001488 => x"03A00000",
001489 => x"0A000000",
001490 => x"EAFFFFF5",
001491 => x"E8FD8070",
001492 => x"07000000",
001493 => x"F0000000",
001494 => x"FFFF0200",
001495 => x"FFFF0218",
001496 => x"E3520007",
001497 => x"E92D45F0",
001498 => x"E1A0C001",
001499 => x"E1A04002",
001500 => x"E1A0A000",
001501 => x"E1A0E000",
001502 => x"83A02000",
001503 => x"8A00001E",
001504 => x"E2443001",
001505 => x"E3530006",
001506 => x"979FF103",
001507 => x"EA000140",
001508 => x"000117E4",
001509 => x"000117DC",
001510 => x"000117D4",
001511 => x"000117CC",
001512 => x"000117C4",
001513 => x"000117BC",
001514 => x"000117AC",
001515 => x"E4D13001",
001516 => x"E1A0E000",
001517 => x"E4CE3001",
001518 => x"E1A0C001",
001519 => x"E4DC3001",
001520 => x"E4CE3001",
001521 => x"E4DC3001",
001522 => x"E4CE3001",
001523 => x"E4DC3001",
001524 => x"E4CE3001",
001525 => x"E4DC3001",
001526 => x"E4CE3001",
001527 => x"E4DC3001",
001528 => x"E4CE3001",
001529 => x"E5DC3000",
001530 => x"E5CE3000",
001531 => x"EA000128",
001532 => x"E7D23001",
001533 => x"E7C2300A",
001534 => x"E2822001",
001535 => x"E08AE002",
001536 => x"E31E0003",
001537 => x"1AFFFFF9",
001538 => x"E0811002",
001539 => x"E2013003",
001540 => x"E0626004",
001541 => x"E3530003",
001542 => x"979FF103",
001543 => x"EA00011B",
001544 => x"00011830",
001545 => x"00011900",
001546 => x"00011A10",
001547 => x"00011B20",
001548 => x"E1A02126",
001549 => x"E3A0C000",
001550 => x"EA000003",
001551 => x"E79C3001",
001552 => x"E2422001",
001553 => x"E78C300E",
001554 => x"E28CC004",
001555 => x"E3120007",
001556 => x"1AFFFFF9",
001557 => x"E08E500C",
001558 => x"E081100C",
001559 => x"E1A021A2",
001560 => x"E1A0E005",
001561 => x"E1A0C001",
001562 => x"E1A04002",
001563 => x"EA00000F",
001564 => x"E51C3020",
001565 => x"E50E3020",
001566 => x"E51C301C",
001567 => x"E50E301C",
001568 => x"E51C3018",
001569 => x"E50E3018",
001570 => x"E51C3014",
001571 => x"E50E3014",
001572 => x"E51C3010",
001573 => x"E50E3010",
001574 => x"E51C300C",
001575 => x"E50E300C",
001576 => x"E51C3008",
001577 => x"E50E3008",
001578 => x"E51C3004",
001579 => x"E50E3004",
001580 => x"E2444001",
001581 => x"E3740001",
001582 => x"E28EE020",
001583 => x"E28CC020",
001584 => x"1AFFFFEA",
001585 => x"E2063003",
001586 => x"E1A02282",
001587 => x"E2433001",
001588 => x"E085C002",
001589 => x"E0811002",
001590 => x"E3530006",
001591 => x"979FF103",
001592 => x"EA0000EB",
001593 => x"00011C84",
001594 => x"00011C7C",
001595 => x"00011C74",
001596 => x"00011C6C",
001597 => x"00011C64",
001598 => x"00011C5C",
001599 => x"00011C54",
001600 => x"E3C10003",
001601 => x"E5904000",
001602 => x"E3CE1003",
001603 => x"E1A0C126",
001604 => x"E1A02001",
001605 => x"EA000003",
001606 => x"E7954003",
001607 => x"E18E3C04",
001608 => x"E5023004",
001609 => x"E24CC001",
001610 => x"E2822004",
001611 => x"E31C0007",
001612 => x"E2615000",
001613 => x"E1A0E424",
001614 => x"E0803002",
001615 => x"1AFFFFF5",
001616 => x"E0613000",
001617 => x"E0837002",
001618 => x"E1A001AC",
001619 => x"E2428004",
001620 => x"E1A0E008",
001621 => x"E1A0C007",
001622 => x"E1A05000",
001623 => x"EA00001F",
001624 => x"E51C2020",
001625 => x"E1A03C02",
001626 => x"E1833424",
001627 => x"E50E3020",
001628 => x"E51C101C",
001629 => x"E1A03C01",
001630 => x"E1833422",
001631 => x"E50E301C",
001632 => x"E51C2018",
001633 => x"E1A03C02",
001634 => x"E1833421",
001635 => x"E50E3018",
001636 => x"E51C1014",
001637 => x"E1A03C01",
001638 => x"E1833422",
001639 => x"E50E3014",
001640 => x"E51C2010",
001641 => x"E1A03C02",
001642 => x"E1833421",
001643 => x"E50E3010",
001644 => x"E51C100C",
001645 => x"E1A03C01",
001646 => x"E1833422",
001647 => x"E50E300C",
001648 => x"E51C2008",
001649 => x"E1A03C02",
001650 => x"E1833421",
001651 => x"E50E3008",
001652 => x"E51C4004",
001653 => x"E1A03C04",
001654 => x"E1833422",
001655 => x"E50E3004",
001656 => x"E2455001",
001657 => x"E3750001",
001658 => x"E28EE020",
001659 => x"E28CC020",
001660 => x"1AFFFFDA",
001661 => x"E1A03280",
001662 => x"E2062003",
001663 => x"E0871003",
001664 => x"E2422001",
001665 => x"E088C003",
001666 => x"E2411003",
001667 => x"EA000086",
001668 => x"E3C10003",
001669 => x"E5904000",
001670 => x"E3CE1003",
001671 => x"E1A0C126",
001672 => x"E1A02001",
001673 => x"EA000003",
001674 => x"E7954003",
001675 => x"E18E3804",
001676 => x"E5023004",
001677 => x"E24CC001",
001678 => x"E2822004",
001679 => x"E31C0007",
001680 => x"E2615000",
001681 => x"E1A0E824",
001682 => x"E0803002",
001683 => x"1AFFFFF5",
001684 => x"E0613000",
001685 => x"E0837002",
001686 => x"E1A001AC",
001687 => x"E2428004",
001688 => x"E1A0E008",
001689 => x"E1A0C007",
001690 => x"E1A05000",
001691 => x"EA00001F",
001692 => x"E51C2020",
001693 => x"E1A03802",
001694 => x"E1833824",
001695 => x"E50E3020",
001696 => x"E51C101C",
001697 => x"E1A03801",
001698 => x"E1833822",
001699 => x"E50E301C",
001700 => x"E51C2018",
001701 => x"E1A03802",
001702 => x"E1833821",
001703 => x"E50E3018",
001704 => x"E51C1014",
001705 => x"E1A03801",
001706 => x"E1833822",
001707 => x"E50E3014",
001708 => x"E51C2010",
001709 => x"E1A03802",
001710 => x"E1833821",
001711 => x"E50E3010",
001712 => x"E51C100C",
001713 => x"E1A03801",
001714 => x"E1833822",
001715 => x"E50E300C",
001716 => x"E51C2008",
001717 => x"E1A03802",
001718 => x"E1833821",
001719 => x"E50E3008",
001720 => x"E51C4004",
001721 => x"E1A03804",
001722 => x"E1833822",
001723 => x"E50E3004",
001724 => x"E2455001",
001725 => x"E3750001",
001726 => x"E28EE020",
001727 => x"E28CC020",
001728 => x"1AFFFFDA",
001729 => x"E1A03280",
001730 => x"E2062003",
001731 => x"E0871003",
001732 => x"E2422001",
001733 => x"E088C003",
001734 => x"E2411002",
001735 => x"EA000042",
001736 => x"E3C10003",
001737 => x"E5904000",
001738 => x"E3CE1003",
001739 => x"E1A0C126",
001740 => x"E1A02001",
001741 => x"EA000003",
001742 => x"E7954003",
001743 => x"E18E3404",
001744 => x"E5023004",
001745 => x"E24CC001",
001746 => x"E2822004",
001747 => x"E31C0007",
001748 => x"E2615000",
001749 => x"E1A0EC24",
001750 => x"E0803002",
001751 => x"1AFFFFF5",
001752 => x"E0613000",
001753 => x"E0837002",
001754 => x"E1A001AC",
001755 => x"E2428004",
001756 => x"E1A0E008",
001757 => x"E1A0C007",
001758 => x"E1A05000",
001759 => x"EA00001F",
001760 => x"E51C2020",
001761 => x"E1A03402",
001762 => x"E1833C24",
001763 => x"E50E3020",
001764 => x"E51C101C",
001765 => x"E1A03401",
001766 => x"E1833C22",
001767 => x"E50E301C",
001768 => x"E51C2018",
001769 => x"E1A03402",
001770 => x"E1833C21",
001771 => x"E50E3018",
001772 => x"E51C1014",
001773 => x"E1A03401",
001774 => x"E1833C22",
001775 => x"E50E3014",
001776 => x"E51C2010",
001777 => x"E1A03402",
001778 => x"E1833C21",
001779 => x"E50E3010",
001780 => x"E51C100C",
001781 => x"E1A03401",
001782 => x"E1833C22",
001783 => x"E50E300C",
001784 => x"E51C2008",
001785 => x"E1A03402",
001786 => x"E1833C21",
001787 => x"E50E3008",
001788 => x"E51C4004",
001789 => x"E1A03404",
001790 => x"E1833C22",
001791 => x"E50E3004",
001792 => x"E2455001",
001793 => x"E3750001",
001794 => x"E28EE020",
001795 => x"E28CC020",
001796 => x"1AFFFFDA",
001797 => x"E1A03280",
001798 => x"E2062003",
001799 => x"E0871003",
001800 => x"E2422001",
001801 => x"E088C003",
001802 => x"E2411001",
001803 => x"E3520006",
001804 => x"979FF102",
001805 => x"EA000016",
001806 => x"00011C84",
001807 => x"00011C7C",
001808 => x"00011C74",
001809 => x"00011C6C",
001810 => x"00011C64",
001811 => x"00011C5C",
001812 => x"00011C54",
001813 => x"E4D13001",
001814 => x"E4CC3001",
001815 => x"E4D13001",
001816 => x"E4CC3001",
001817 => x"E4D13001",
001818 => x"E4CC3001",
001819 => x"E4D13001",
001820 => x"E4CC3001",
001821 => x"E4D13001",
001822 => x"E4CC3001",
001823 => x"E4D13001",
001824 => x"E4CC3001",
001825 => x"E5D13000",
001826 => x"E5CC3000",
001827 => x"EA000000",
001828 => x"E8BD85F0",
001829 => x"E1A0000A",
001830 => x"E8BD85F0",
001831 => x"00001021",
001832 => x"20423063",
001833 => x"408450A5",
001834 => x"60C670E7",
001835 => x"81089129",
001836 => x"A14AB16B",
001837 => x"C18CD1AD",
001838 => x"E1CEF1EF",
001839 => x"12310210",
001840 => x"32732252",
001841 => x"52B54294",
001842 => x"72F762D6",
001843 => x"93398318",
001844 => x"B37BA35A",
001845 => x"D3BDC39C",
001846 => x"F3FFE3DE",
001847 => x"24623443",
001848 => x"04201401",
001849 => x"64E674C7",
001850 => x"44A45485",
001851 => x"A56AB54B",
001852 => x"85289509",
001853 => x"E5EEF5CF",
001854 => x"C5ACD58D",
001855 => x"36532672",
001856 => x"16110630",
001857 => x"76D766F6",
001858 => x"569546B4",
001859 => x"B75BA77A",
001860 => x"97198738",
001861 => x"F7DFE7FE",
001862 => x"D79DC7BC",
001863 => x"48C458E5",
001864 => x"688678A7",
001865 => x"08401861",
001866 => x"28023823",
001867 => x"C9CCD9ED",
001868 => x"E98EF9AF",
001869 => x"89489969",
001870 => x"A90AB92B",
001871 => x"5AF54AD4",
001872 => x"7AB76A96",
001873 => x"1A710A50",
001874 => x"3A332A12",
001875 => x"DBFDCBDC",
001876 => x"FBBFEB9E",
001877 => x"9B798B58",
001878 => x"BB3BAB1A",
001879 => x"6CA67C87",
001880 => x"4CE45CC5",
001881 => x"2C223C03",
001882 => x"0C601C41",
001883 => x"EDAEFD8F",
001884 => x"CDECDDCD",
001885 => x"AD2ABD0B",
001886 => x"8D689D49",
001887 => x"7E976EB6",
001888 => x"5ED54EF4",
001889 => x"3E132E32",
001890 => x"1E510E70",
001891 => x"FF9FEFBE",
001892 => x"DFDDCFFC",
001893 => x"BF1BAF3A",
001894 => x"9F598F78",
001895 => x"918881A9",
001896 => x"B1CAA1EB",
001897 => x"D10CC12D",
001898 => x"F14EE16F",
001899 => x"108000A1",
001900 => x"30C220E3",
001901 => x"50044025",
001902 => x"70466067",
001903 => x"83B99398",
001904 => x"A3FBB3DA",
001905 => x"C33DD31C",
001906 => x"E37FF35E",
001907 => x"02B11290",
001908 => x"22F332D2",
001909 => x"42355214",
001910 => x"62777256",
001911 => x"B5EAA5CB",
001912 => x"95A88589",
001913 => x"F56EE54F",
001914 => x"D52CC50D",
001915 => x"34E224C3",
001916 => x"14A00481",
001917 => x"74666447",
001918 => x"54244405",
001919 => x"A7DBB7FA",
001920 => x"879997B8",
001921 => x"E75FF77E",
001922 => x"C71DD73C",
001923 => x"26D336F2",
001924 => x"069116B0",
001925 => x"66577676",
001926 => x"46155634",
001927 => x"D94CC96D",
001928 => x"F90EE92F",
001929 => x"99C889E9",
001930 => x"B98AA9AB",
001931 => x"58444865",
001932 => x"78066827",
001933 => x"18C008E1",
001934 => x"388228A3",
001935 => x"CB7DDB5C",
001936 => x"EB3FFB1E",
001937 => x"8BF99BD8",
001938 => x"ABBBBB9A",
001939 => x"4A755A54",
001940 => x"6A377A16",
001941 => x"0AF11AD0",
001942 => x"2AB33A92",
001943 => x"FD2EED0F",
001944 => x"DD6CCD4D",
001945 => x"BDAAAD8B",
001946 => x"9DE88DC9",
001947 => x"7C266C07",
001948 => x"5C644C45",
001949 => x"3CA22C83",
001950 => x"1CE00CC1",
001951 => x"EF1FFF3E",
001952 => x"CF5DDF7C",
001953 => x"AF9BBFBA",
001954 => x"8FD99FF8",
001955 => x"6E177E36",
001956 => x"4E555E74",
001957 => x"2E933EB2",
001958 => x"0ED11EF0",
001959 => x"25632000",
001960 => x"20000000",
001961 => x"436F6D6D",
001962 => x"616E6473",
001963 => x"0A000000",
001964 => x"6C000000",
001965 => x"3A204C6F",
001966 => x"61642065",
001967 => x"6C662066",
001968 => x"696C650A",
001969 => x"00000000",
001970 => x"62203C61",
001971 => x"64647265",
001972 => x"73733E00",
001973 => x"3A204C6F",
001974 => x"61642062",
001975 => x"696E6172",
001976 => x"79206669",
001977 => x"6C652074",
001978 => x"6F203C61",
001979 => x"64647265",
001980 => x"73733E0A",
001981 => x"00000000",
001982 => x"64203C73",
001983 => x"74617274",
001984 => x"20616464",
001985 => x"72657373",
001986 => x"3E203C6E",
001987 => x"756D2062",
001988 => x"79746573",
001989 => x"3E203A20",
001990 => x"44756D70",
001991 => x"206D656D",
001992 => x"0A000000",
001993 => x"68000000",
001994 => x"3A205072",
001995 => x"696E7420",
001996 => x"68656C70",
001997 => x"206D6573",
001998 => x"73616765",
001999 => x"0A000000",
002000 => x"6A203C61",
002001 => x"64647265",
002002 => x"73733E00",
002003 => x"3A204578",
002004 => x"65637574",
002005 => x"65206C6F",
002006 => x"61646564",
002007 => x"20656C66",
002008 => x"2C206A75",
002009 => x"6D70696E",
002010 => x"6720746F",
002011 => x"203C6164",
002012 => x"64726573",
002013 => x"733E0A00",
002014 => x"70203C61",
002015 => x"64647265",
002016 => x"73733E00",
002017 => x"3A205072",
002018 => x"696E7420",
002019 => x"61736369",
002020 => x"69206D65",
002021 => x"6D20756E",
002022 => x"74696C20",
002023 => x"66697273",
002024 => x"7420300A",
002025 => x"00000000",
002026 => x"72203C61",
002027 => x"64647265",
002028 => x"73733E00",
002029 => x"3A205265",
002030 => x"6164206D",
002031 => x"656D0A00",
002032 => x"73000000",
002033 => x"3A20436F",
002034 => x"72652073",
002035 => x"74617475",
002036 => x"730A0000",
002037 => x"77203C61",
002038 => x"64647265",
002039 => x"73733E20",
002040 => x"3C76616C",
002041 => x"75653E00",
002042 => x"3A205772",
002043 => x"69746520",
002044 => x"6D656D0A",
002045 => x"00000000",
002046 => x"61646472",
002047 => x"6573733A",
002048 => x"20257820",
002049 => x"0A000000",
002050 => x"6D656D20",
002051 => x"30782530",
002052 => x"3878203D",
002053 => x"20307825",
002054 => x"3038780A",
002055 => x"00000000",
002056 => x"25730A00",
002057 => x"53656E64",
002058 => x"2066696C",
002059 => x"6520772F",
002060 => x"20314B20",
002061 => x"586D6F64",
002062 => x"656D2070",
002063 => x"726F746F",
002064 => x"636F6C20",
002065 => x"66726F6D",
002066 => x"20746572",
002067 => x"6D696E61",
002068 => x"6C20656D",
002069 => x"756C6174",
002070 => x"6F72206E",
002071 => x"6F772E2E",
002072 => x"2E000000",
002073 => x"586D6F64",
002074 => x"656D2065",
002075 => x"72726F72",
002076 => x"2066696C",
002077 => x"65207369",
002078 => x"7A652030",
002079 => x"78257820",
002080 => x"0A000000",
002081 => x"0A656C66",
002082 => x"2073706C",
002083 => x"69740A00",
002084 => x"6A203078",
002085 => x"25303878",
002086 => x"0A000000",
002087 => x"64617461",
002088 => x"3A202578",
002089 => x"202D6E00",
002090 => x"496E7661",
002091 => x"6C696420",
002092 => x"636F6D6D",
002093 => x"616E6400",
002094 => x"2563416D",
002095 => x"62657220",
002096 => x"426F6F74",
002097 => x"204C6F61",
002098 => x"64657220",
002099 => x"77697468",
002100 => x"20444530",
002101 => x"2D4E414E",
002102 => x"4F203332",
002103 => x"4D422073",
002104 => x"7570706F",
002105 => x"72747625",
002106 => x"730A0000",
002107 => x"32303135",
002108 => x"2D30392D",
002109 => x"31370000",
002110 => x"52656164",
002111 => x"790A3E20",
002112 => x"00000000",
002113 => x"3E200000",
002114 => x"44656275",
002115 => x"673A2073",
002116 => x"697A6520",
002117 => x"3D202564",
002118 => x"0A000000",
002119 => x"44656275",
002120 => x"673A2065",
002121 => x"6C664865",
002122 => x"61646572",
002123 => x"2D3E655F",
002124 => x"6D616368",
002125 => x"696E653D",
002126 => x"20307825",
002127 => x"780A0000",
002128 => x"454C4600",
002129 => x"4552524F",
002130 => x"523A204E",
002131 => x"6F742061",
002132 => x"6E20454C",
002133 => x"46206669",
002134 => x"6C652E0A",
002135 => x"00000000",
002136 => x"4552524F",
002137 => x"523A2045",
002138 => x"4C462066",
002139 => x"696C6520",
002140 => x"6E6F7420",
002141 => x"74617267",
002142 => x"65747469",
002143 => x"6E672063",
002144 => x"6F727265",
002145 => x"63742070",
002146 => x"726F6365",
002147 => x"73736F72",
002148 => x"20747970",
002149 => x"650A0000",
002150 => x"44656275",
002151 => x"673A2065",
002152 => x"6C664865",
002153 => x"61646572",
002154 => x"2D3E655F",
002155 => x"70686E75",
002156 => x"6D3D3078",
002157 => x"25780A00",
002158 => x"44656275",
002159 => x"673A2050",
002160 => x"726F6772",
002161 => x"616D204C",
002162 => x"656E6774",
002163 => x"683D3078",
002164 => x"25780A00",
002165 => x"286E756C",
002166 => x"6C290000",
others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;