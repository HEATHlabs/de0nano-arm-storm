-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
--				MEM_SIZE      : natural := 1024;  -- memory cells
--				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				MEM_SIZE      : natural := 2048;  -- memory cells
				LOG2_MEM_SIZE : natural := 11;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
000000 => x"EA000006",
000001 => x"EA00047B",
000002 => x"EA00047A",
000003 => x"EA000479",
000004 => x"EA000478",
000005 => x"EA000477",
000006 => x"EA000476",
000007 => x"EA000475",
000008 => x"E59F0168",
000009 => x"E10F1000",
000010 => x"E3C1107F",
000011 => x"E38110DF",
000012 => x"E129F001",
000013 => x"E1A0D000",
000014 => x"E3A00000",
000015 => x"E1A01000",
000016 => x"E1A02000",
000017 => x"E1A0B000",
000018 => x"E1A07000",
000019 => x"E59FA140",
000020 => x"E1A0E00F",
000021 => x"E1A0F00A",
000022 => x"E3A00003",
000023 => x"E13FF000",
000024 => x"E59FD098",
000025 => x"EB0001D6",
000026 => x"E59F1118",
000027 => x"E59F20B8",
000028 => x"E59F30B8",
000029 => x"E1520003",
000030 => x"0A000002",
000031 => x"E4924004",
000032 => x"E4814004",
000033 => x"EAFFFFFA",
000034 => x"E59F20FC",
000035 => x"E3A03000",
000036 => x"E3A04028",
000037 => x"E4823004",
000038 => x"E2544001",
000039 => x"1AFFFFFC",
000040 => x"E1A04000",
000041 => x"E38443C3",
000042 => x"E3A00000",
000043 => x"E1A0F004",
000044 => x"E92D4000",
000045 => x"E92D1FFF",
000046 => x"E3A04000",
000047 => x"E1A0500D",
000048 => x"E1A0600E",
000049 => x"E59F00CC",
000050 => x"E1A01004",
000051 => x"E4952004",
000052 => x"EB00042D",
000053 => x"E354000D",
000054 => x"12844001",
000055 => x"1AFFFFF8",
000056 => x"E59F00B4",
000057 => x"E1A0100D",
000058 => x"EB000427",
000059 => x"E59F00AC",
000060 => x"E2461004",
000061 => x"EB000424",
000062 => x"E8BD1FFF",
000063 => x"E8FD8000",
000064 => x"007FFFF8",
000065 => x"F0000020",
000066 => x"72253264",
000067 => x"20202530",
000068 => x"38780A00",
000069 => x"73702020",
000070 => x"20253038",
000071 => x"780A0070",
000072 => x"63202020",
000073 => x"25303878",
000074 => x"0A000000",
000075 => x"00010134",
000076 => x"00010184",
000077 => x"00000005",
000078 => x"54410001",
000079 => x"00000001",
000080 => x"00001000",
000081 => x"00000000",
000082 => x"00000004",
000083 => x"54410002",
000084 => x"00800000",
000085 => x"00000000",
000086 => x"00000005",
000087 => x"54410004",
000088 => x"00000001",
000089 => x"000000D0",
000090 => x"00001E00",
000091 => x"00000004",
000092 => x"54410005",
000093 => x"02700000",
000094 => x"00034000",
000095 => x"00000000",
000096 => x"00000000",
000097 => x"00000000",
000098 => x"0007C000",
000099 => x"03F01000",
000100 => x"00002100",
000101 => x"000107C4",
000102 => x"00010108",
000103 => x"00010114",
000104 => x"0001011F",
000105 => x"E1A0C002",
000106 => x"E3A02000",
000107 => x"E58C2000",
000108 => x"E92D40F0",
000109 => x"E0800001",
000110 => x"E1A06003",
000111 => x"E1A04002",
000112 => x"E1A05001",
000113 => x"E5D02000",
000114 => x"E2423030",
000115 => x"E3530009",
000116 => x"E242E041",
000117 => x"E3A07000",
000118 => x"8A000006",
000119 => x"E59C3000",
000120 => x"E1A03203",
000121 => x"E58C3000",
000122 => x"E5D02000",
000123 => x"E0833002",
000124 => x"E2433030",
000125 => x"EA000009",
000126 => x"E35E0005",
000127 => x"E2423061",
000128 => x"E3A07000",
000129 => x"8A000007",
000130 => x"E59C3000",
000131 => x"E1A03203",
000132 => x"E58C3000",
000133 => x"E5D02000",
000134 => x"E0833002",
000135 => x"E2433037",
000136 => x"E58C3000",
000137 => x"EA00000B",
000138 => x"E3530005",
000139 => x"E3A07000",
000140 => x"85864000",
000141 => x"83A07001",
000142 => x"8A000006",
000143 => x"E59C3000",
000144 => x"E1A03203",
000145 => x"E58C3000",
000146 => x"E5D02000",
000147 => x"E0833002",
000148 => x"E2433057",
000149 => x"EAFFFFF1",
000150 => x"E2853001",
000151 => x"E3540008",
000152 => x"E2800001",
000153 => x"E1A05003",
000154 => x"05864000",
000155 => x"0A000002",
000156 => x"E3570000",
000157 => x"E2844001",
000158 => x"0AFFFFD1",
000159 => x"E2810001",
000160 => x"E1530000",
000161 => x"D3A00000",
000162 => x"C3A00001",
000163 => x"E8BD80F0",
000164 => x"E92D4070",
000165 => x"E24DD004",
000166 => x"E1A06002",
000167 => x"E1A0300D",
000168 => x"E1A02001",
000169 => x"E3A01002",
000170 => x"E1A04000",
000171 => x"EBFFFFBC",
000172 => x"E2501000",
000173 => x"E1A0500D",
000174 => x"E1A02006",
000175 => x"E1A00004",
000176 => x"E1A0300D",
000177 => x"0A000003",
000178 => x"E59D1000",
000179 => x"E2811003",
000180 => x"EBFFFFB3",
000181 => x"E1A01000",
000182 => x"E1A00001",
000183 => x"E28DD004",
000184 => x"E8BD8070",
000185 => x"E92D4010",
000186 => x"E1A04000",
000187 => x"EA000000",
000188 => x"EB0003A5",
000189 => x"E2544001",
000190 => x"E59F0004",
000191 => x"2AFFFFFB",
000192 => x"E8BD8010",
000193 => x"00011DB4",
000194 => x"E52DE004",
000195 => x"E59F00CC",
000196 => x"EB00039D",
000197 => x"E59F00C8",
000198 => x"EB00039B",
000199 => x"E3A0001D",
000200 => x"EBFFFFEF",
000201 => x"E59F00BC",
000202 => x"EB000397",
000203 => x"E59F00B8",
000204 => x"EB000395",
000205 => x"E3A00013",
000206 => x"EBFFFFE9",
000207 => x"E59F00AC",
000208 => x"EB000391",
000209 => x"E59F00A8",
000210 => x"EB00038F",
000211 => x"E59F00A4",
000212 => x"EB00038D",
000213 => x"E3A0001D",
000214 => x"EBFFFFE1",
000215 => x"E59F0098",
000216 => x"EB000389",
000217 => x"E59F0094",
000218 => x"EB000387",
000219 => x"E3A00013",
000220 => x"EBFFFFDB",
000221 => x"E59F0088",
000222 => x"EB000383",
000223 => x"E59F0084",
000224 => x"EB000381",
000225 => x"E3A00013",
000226 => x"EBFFFFD5",
000227 => x"E59F0078",
000228 => x"EB00037D",
000229 => x"E59F0074",
000230 => x"EB00037B",
000231 => x"E3A00013",
000232 => x"EBFFFFCF",
000233 => x"E59F0068",
000234 => x"EB000377",
000235 => x"E59F0064",
000236 => x"EB000375",
000237 => x"E3A0001D",
000238 => x"EBFFFFC9",
000239 => x"E59F0058",
000240 => x"EB000371",
000241 => x"E59F0054",
000242 => x"EB00036F",
000243 => x"E3A0000B",
000244 => x"EBFFFFC3",
000245 => x"E59F0048",
000246 => x"E49DE004",
000247 => x"EA00036A",
000248 => x"00011DB8",
000249 => x"00011DC4",
000250 => x"00011DC8",
000251 => x"00011DDC",
000252 => x"00011DE8",
000253 => x"00011E0C",
000254 => x"00011E38",
000255 => x"00011E3C",
000256 => x"00011E54",
000257 => x"00011E60",
000258 => x"00011E8C",
000259 => x"00011E98",
000260 => x"00011EBC",
000261 => x"00011EC8",
000262 => x"00011ED4",
000263 => x"00011ED8",
000264 => x"00011EE8",
000265 => x"00011EFC",
000266 => x"E1A01000",
000267 => x"E5912000",
000268 => x"E59F0000",
000269 => x"EA000354",
000270 => x"00011F0C",
000271 => x"E2400001",
000272 => x"E92D4010",
000273 => x"E1A04001",
000274 => x"E3500004",
000275 => x"979FF100",
000276 => x"EA000039",
000277 => x"00010468",
000278 => x"000104A8",
000279 => x"000104BC",
000280 => x"000104E8",
000281 => x"0001050C",
000282 => x"E59F10EC",
000283 => x"E59F00EC",
000284 => x"EB000345",
000285 => x"E3A01602",
000286 => x"E3A00505",
000287 => x"EB000153",
000288 => x"E3500602",
000289 => x"E1A04000",
000290 => x"81A01000",
000291 => x"8A000027",
000292 => x"E59F00CC",
000293 => x"EB00033C",
000294 => x"E1A01004",
000295 => x"E3A00505",
000296 => x"E8BD4010",
000297 => x"EA0001EE",
000298 => x"EBFFFF96",
000299 => x"EBFFFEFF",
000300 => x"E3A00010",
000301 => x"EBFFFF8A",
000302 => x"EA000008",
000303 => x"E3A01702",
000304 => x"E59F00A0",
000305 => x"EB000330",
000306 => x"E3A00010",
000307 => x"EBFFFF84",
000308 => x"E59F0094",
000309 => x"EB00032C",
000310 => x"E3A00702",
000311 => x"EBFFFEE1",
000312 => x"E8BD4010",
000313 => x"EA000346",
000314 => x"E3A01901",
000315 => x"E59F0074",
000316 => x"EB000325",
000317 => x"E3A00010",
000318 => x"EBFFFF79",
000319 => x"E59F0068",
000320 => x"EB000321",
000321 => x"E3A00901",
000322 => x"EAFFFFF3",
000323 => x"E59F1048",
000324 => x"E59F0048",
000325 => x"EB00031C",
000326 => x"E1A00004",
000327 => x"E3A01602",
000328 => x"EB00012A",
000329 => x"E3500602",
000330 => x"98BD8010",
000331 => x"E1A01000",
000332 => x"E59F0038",
000333 => x"E8BD4010",
000334 => x"EA000313",
000335 => x"E59F0024",
000336 => x"EB000311",
000337 => x"E3A00010",
000338 => x"EBFFFF65",
000339 => x"E59F0018",
000340 => x"EB00030D",
000341 => x"E1A00004",
000342 => x"EAFFFFDF",
000343 => x"00011F28",
000344 => x"00011F24",
000345 => x"00011F88",
000346 => x"00011F94",
000347 => x"00011F84",
000348 => x"00011F68",
000349 => x"E92D4010",
000350 => x"E59F3238",
000351 => x"E5D0C001",
000352 => x"E1A0E000",
000353 => x"E893000F",
000354 => x"E24DD020",
000355 => x"E35C0000",
000356 => x"E1A0400D",
000357 => x"E88D000F",
000358 => x"0A000084",
000359 => x"E35C000D",
000360 => x"1A000011",
000361 => x"E5DE0000",
000362 => x"E350006C",
000363 => x"0A000005",
000364 => x"E3500073",
000365 => x"0A000006",
000366 => x"E3500068",
000367 => x"1A00000C",
000368 => x"EBFFFF50",
000369 => x"EA000079",
000370 => x"E3A00001",
000371 => x"E3A01000",
000372 => x"EA000034",
000373 => x"EBFFFEB5",
000374 => x"E3A00010",
000375 => x"EBFFFF40",
000376 => x"E59F01D4",
000377 => x"EB0002E8",
000378 => x"EA000070",
000379 => x"E35C0020",
000380 => x"0A000002",
000381 => x"E59F01C4",
000382 => x"E1A0100D",
000383 => x"EA00006A",
000384 => x"E5DE3000",
000385 => x"E353006A",
000386 => x"0A00001D",
000387 => x"8A000004",
000388 => x"E3530062",
000389 => x"0A00004D",
000390 => x"E3530064",
000391 => x"1A000060",
000392 => x"EA000006",
000393 => x"E3530072",
000394 => x"0A000040",
000395 => x"E3530077",
000396 => x"0A00004F",
000397 => x"E3530070",
000398 => x"1A000059",
000399 => x"EA00001B",
000400 => x"E1A0000E",
000401 => x"E28D1010",
000402 => x"E28D2014",
000403 => x"EBFFFF0F",
000404 => x"E3500000",
000405 => x"159D4010",
000406 => x"1A000001",
000407 => x"EA000053",
000408 => x"EBFFFF70",
000409 => x"E59D3010",
000410 => x"E59D2014",
000411 => x"E0833002",
000412 => x"E1540003",
000413 => x"E1A00004",
000414 => x"E2844004",
000415 => x"3AFFFFF7",
000416 => x"EA00004A",
000417 => x"E1A0000E",
000418 => x"E3A01002",
000419 => x"E28D2010",
000420 => x"E28D3018",
000421 => x"EBFFFEC2",
000422 => x"E3500000",
000423 => x"0A000043",
000424 => x"E3A00000",
000425 => x"E59D1010",
000426 => x"EBFFFF63",
000427 => x"EA00003F",
000428 => x"E1A0000E",
000429 => x"E3A01002",
000430 => x"E28D2010",
000431 => x"E28D3018",
000432 => x"EBFFFEB7",
000433 => x"E3500000",
000434 => x"0A000038",
000435 => x"E3A03000",
000436 => x"E58D3018",
000437 => x"E59D3010",
000438 => x"E4D34001",
000439 => x"E58D3010",
000440 => x"EA00000B",
000441 => x"E3540000",
000442 => x"0A000003",
000443 => x"EB0002C8",
000444 => x"E354000D",
000445 => x"E59F00C0",
000446 => x"0B0002A3",
000447 => x"E59D2010",
000448 => x"E59D3018",
000449 => x"E4D24001",
000450 => x"E2833001",
000451 => x"E58D2010",
000452 => x"E58D3018",
000453 => x"E3140080",
000454 => x"E1A00004",
000455 => x"1A000023",
000456 => x"E59D3018",
000457 => x"E3530A01",
000458 => x"3AFFFFED",
000459 => x"EA00001F",
000460 => x"E1A0000E",
000461 => x"E3A01002",
000462 => x"E28D2010",
000463 => x"E28D3018",
000464 => x"EBFFFE97",
000465 => x"E3500000",
000466 => x"0A000018",
000467 => x"EA000011",
000468 => x"E1A0000E",
000469 => x"E3A01002",
000470 => x"E28D2010",
000471 => x"E28D3018",
000472 => x"EBFFFE8F",
000473 => x"E3500000",
000474 => x"13A00005",
000475 => x"1AFFFFCC",
000476 => x"EA00000E",
000477 => x"E1A0000E",
000478 => x"E28D1010",
000479 => x"E28D201C",
000480 => x"EBFFFEC2",
000481 => x"E3500000",
000482 => x"0A000008",
000483 => x"E59D201C",
000484 => x"E59D3010",
000485 => x"E5832000",
000486 => x"E59D0010",
000487 => x"EBFFFF21",
000488 => x"EA000002",
000489 => x"E59F0014",
000490 => x"E1A0100D",
000491 => x"EB000276",
000492 => x"E28DD020",
000493 => x"E8BD8010",
000494 => x"00011FA0",
000495 => x"00011F84",
000496 => x"00011F24",
000497 => x"E92D41F0",
000498 => x"E3A0100C",
000499 => x"E24DD028",
000500 => x"E59F2170",
000501 => x"E59F0170",
000502 => x"EB00026B",
000503 => x"EBFFFEC9",
000504 => x"E59F0168",
000505 => x"EB000268",
000506 => x"E3A06000",
000507 => x"E1A07006",
000508 => x"E1A08006",
000509 => x"EA000001",
000510 => x"E1A06008",
000511 => x"E3A07000",
000512 => x"E3A00FFA",
000513 => x"EB00028A",
000514 => x"E2504000",
000515 => x"BAFFFFFB",
000516 => x"E354001B",
000517 => x"0A00001C",
000518 => x"E3570001",
000519 => x"0354005B",
000520 => x"13A05000",
000521 => x"03A05001",
000522 => x"03A07002",
000523 => x"0A00001D",
000524 => x"E3570002",
000525 => x"1A000038",
000526 => x"E3540041",
000527 => x"01A04005",
000528 => x"11A07005",
000529 => x"1AFFFFED",
000530 => x"EA000000",
000531 => x"EB000270",
000532 => x"E1540006",
000533 => x"E3A00008",
000534 => x"E2844001",
000535 => x"BAFFFFFA",
000536 => x"E3A04000",
000537 => x"EA000005",
000538 => x"E28D3014",
000539 => x"E7D42003",
000540 => x"E1A00002",
000541 => x"E7C4200D",
000542 => x"EB000265",
000543 => x"E2844001",
000544 => x"E1540008",
000545 => x"BAFFFFF7",
000546 => x"EAFFFFDA",
000547 => x"E3A07001",
000548 => x"EA000004",
000549 => x"E28D2028",
000550 => x"E0823006",
000551 => x"E5434028",
000552 => x"E2866001",
000553 => x"E3A07000",
000554 => x"E3560012",
000555 => x"D3A03000",
000556 => x"C3A03001",
000557 => x"E354000D",
000558 => x"03833001",
000559 => x"E3530000",
000560 => x"0AFFFFCE",
000561 => x"E3560001",
000562 => x"DA000007",
000563 => x"E3A01000",
000564 => x"E7D1200D",
000565 => x"E28D3014",
000566 => x"E7C12003",
000567 => x"E2811001",
000568 => x"E3510014",
000569 => x"1AFFFFF9",
000570 => x"E2468001",
000571 => x"E28D2028",
000572 => x"E0823006",
000573 => x"E3A04000",
000574 => x"E5434028",
000575 => x"E59F0050",
000576 => x"EB000221",
000577 => x"E1A0000D",
000578 => x"EBFFFF19",
000579 => x"E59F0044",
000580 => x"EB00021D",
000581 => x"E1A06004",
000582 => x"EAFFFFB8",
000583 => x"EB00023C",
000584 => x"E3540008",
000585 => x"13A03000",
000586 => x"03A03001",
000587 => x"E3560000",
000588 => x"D3A03000",
000589 => x"E3530000",
000590 => x"12466001",
000591 => x"11A07005",
000592 => x"1AFFFFD8",
000593 => x"EAFFFFD2",
000594 => x"00011FE4",
000595 => x"00011FB0",
000596 => x"00011FF0",
000597 => x"00011F84",
000598 => x"00011FFC",
000599 => x"E92D4010",
000600 => x"E3A0C000",
000601 => x"E1A04000",
000602 => x"E1A0E00C",
000603 => x"E1A00001",
000604 => x"EA00000A",
000605 => x"E7DE3004",
000606 => x"E023342C",
000607 => x"E1A03083",
000608 => x"E0832001",
000609 => x"E7D31001",
000610 => x"E5D23001",
000611 => x"E1833401",
000612 => x"E023340C",
000613 => x"E1A03803",
000614 => x"E28EE001",
000615 => x"E1A0C823",
000616 => x"E15E0000",
000617 => x"E59F1008",
000618 => x"BAFFFFF1",
000619 => x"E1A0000C",
000620 => x"E8BD8010",
000621 => x"00011BB4",
000622 => x"E52DE004",
000623 => x"E3A00F4B",
000624 => x"EB00021B",
000625 => x"E3500000",
000626 => x"AAFFFFFB",
000627 => x"E49DF004",
000628 => x"E92D4FF0",
000629 => x"E3A07000",
000630 => x"E24DDB01",
000631 => x"E24DD008",
000632 => x"E1A0B000",
000633 => x"E1A09001",
000634 => x"E3A0A019",
000635 => x"E3A04043",
000636 => x"E3A08001",
000637 => x"E1A06007",
000638 => x"EA000000",
000639 => x"E3A04015",
000640 => x"E3A05000",
000641 => x"E3540000",
000642 => x"11A00004",
000643 => x"1B000200",
000644 => x"E3A00FFA",
000645 => x"EB000206",
000646 => x"E3500000",
000647 => x"BA000019",
000648 => x"E3500002",
000649 => x"0A000025",
000650 => x"CA000002",
000651 => x"E3500001",
000652 => x"1A000014",
000653 => x"EA000004",
000654 => x"E3500004",
000655 => x"0A000004",
000656 => x"E3500018",
000657 => x"1A00000F",
000658 => x"EA000005",
000659 => x"E3A05080",
000660 => x"EA00001B",
000661 => x"E3A00006",
000662 => x"EB0001ED",
000663 => x"EBFFFFD5",
000664 => x"EA00007B",
000665 => x"E3A00FFA",
000666 => x"EB0001F1",
000667 => x"E3500018",
000668 => x"1A000004",
000669 => x"EBFFFFCF",
000670 => x"E3A00006",
000671 => x"EB0001E4",
000672 => x"E3E06000",
000673 => x"EA000072",
000674 => x"E2855001",
000675 => x"E3550050",
000676 => x"1AFFFFDB",
000677 => x"E3540043",
000678 => x"0AFFFFD7",
000679 => x"EBFFFFC5",
000680 => x"E3A00018",
000681 => x"EB0001DA",
000682 => x"E3A00018",
000683 => x"EB0001D8",
000684 => x"E3A00018",
000685 => x"EB0001D6",
000686 => x"E3E06001",
000687 => x"EA000064",
000688 => x"E3A05B01",
000689 => x"E3540043",
000690 => x"03A07001",
000691 => x"E1A00000",
000692 => x"E3A04000",
000693 => x"E5CD0002",
000694 => x"EA000006",
000695 => x"EB0001D4",
000696 => x"E28D3008",
000697 => x"E3500000",
000698 => x"E2433006",
000699 => x"E2844001",
000700 => x"BA000052",
000701 => x"E7C40003",
000702 => x"E3570000",
000703 => x"13A03004",
000704 => x"03A03003",
000705 => x"E0853003",
000706 => x"E1540003",
000707 => x"E3A00FFA",
000708 => x"BAFFFFF1",
000709 => x"E5DD3004",
000710 => x"E5DD2003",
000711 => x"E1E03003",
000712 => x"E20330FF",
000713 => x"E1520003",
000714 => x"1A000044",
000715 => x"E1520008",
000716 => x"0A000002",
000717 => x"E2483001",
000718 => x"E1520003",
000719 => x"1A00003F",
000720 => x"E3570000",
000721 => x"E28D4008",
000722 => x"E2444006",
000723 => x"01A01007",
000724 => x"02840003",
000725 => x"01A02001",
000726 => x"0A00000D",
000727 => x"E2840003",
000728 => x"E1A01005",
000729 => x"EBFFFF7C",
000730 => x"E0843005",
000731 => x"E5D32004",
000732 => x"E5D33003",
000733 => x"E0822403",
000734 => x"E1A02802",
000735 => x"E1500822",
000736 => x"1A00002E",
000737 => x"EA00000C",
000738 => x"E5503001",
000739 => x"E0813003",
000740 => x"E20310FF",
000741 => x"E1520005",
000742 => x"E2800001",
000743 => x"E2822001",
000744 => x"BAFFFFF8",
000745 => x"E28D2B01",
000746 => x"E2822008",
000747 => x"E0823005",
000748 => x"E5533403",
000749 => x"E1530001",
000750 => x"1A000020",
000751 => x"E5DD3003",
000752 => x"E1530008",
000753 => x"1A00000F",
000754 => x"E0663009",
000755 => x"E1550003",
000756 => x"B1A04005",
000757 => x"A1A04003",
000758 => x"E3540000",
000759 => x"DA000005",
000760 => x"E28D1008",
000761 => x"E08B0006",
000762 => x"E2411003",
000763 => x"E1A02004",
000764 => x"EB0002A0",
000765 => x"E0866004",
000766 => x"E2883001",
000767 => x"E20380FF",
000768 => x"E3A0A019",
000769 => x"EA00000B",
000770 => x"E24AA001",
000771 => x"E35A0000",
000772 => x"CA000008",
000773 => x"EBFFFF67",
000774 => x"E3A00018",
000775 => x"EB00017C",
000776 => x"E3A00018",
000777 => x"EB00017A",
000778 => x"E3A00018",
000779 => x"EB000178",
000780 => x"E3E06002",
000781 => x"EA000006",
000782 => x"E3A00006",
000783 => x"EA000001",
000784 => x"EBFFFF5C",
000785 => x"E3A00015",
000786 => x"EB000171",
000787 => x"E3A04000",
000788 => x"EAFFFF6A",
000789 => x"E1A00006",
000790 => x"E28DD008",
000791 => x"E28DDB01",
000792 => x"E8BD8FF0",
000793 => x"E92D40F0",
000794 => x"E59F1140",
000795 => x"E1A05000",
000796 => x"E3A02003",
000797 => x"E2800001",
000798 => x"EB00026A",
000799 => x"E3500000",
000800 => x"159F012C",
000801 => x"1A000006",
000802 => x"E5D52012",
000803 => x"E5D53013",
000804 => x"E1833402",
000805 => x"E3530028",
000806 => x"01A07000",
000807 => x"0A00003C",
000808 => x"E59F0110",
000809 => x"EB000138",
000810 => x"E3A00001",
000811 => x"E8BD80F0",
000812 => x"E5952020",
000813 => x"E5D5102E",
000814 => x"E5D5302F",
000815 => x"E0852002",
000816 => x"E1833401",
000817 => x"E0242397",
000818 => x"E5943004",
000819 => x"E3530001",
000820 => x"1A000018",
000821 => x"E5943014",
000822 => x"E3530000",
000823 => x"0A00002B",
000824 => x"E594300C",
000825 => x"E3530000",
000826 => x"13A06000",
000827 => x"1A00000E",
000828 => x"EA000026",
000829 => x"E5942010",
000830 => x"E0862002",
000831 => x"E0851002",
000832 => x"E5D13002",
000833 => x"E5D10003",
000834 => x"E7D5C002",
000835 => x"E1A03803",
000836 => x"E5D12001",
000837 => x"E1833C00",
000838 => x"E594E00C",
000839 => x"E183300C",
000840 => x"E1833402",
000841 => x"E78E3006",
000842 => x"E2866004",
000843 => x"E5943014",
000844 => x"E1560003",
000845 => x"3AFFFFEE",
000846 => x"E5943004",
000847 => x"E3530008",
000848 => x"1A000012",
000849 => x"E5943014",
000850 => x"E3530000",
000851 => x"0A00000F",
000852 => x"E594300C",
000853 => x"E3530000",
000854 => x"15941010",
000855 => x"1A000006",
000856 => x"EA00000A",
000857 => x"E594300C",
000858 => x"E0813003",
000859 => x"E0623003",
000860 => x"E3A02000",
000861 => x"E5832000",
000862 => x"E2811004",
000863 => x"E2842010",
000864 => x"E892000C",
000865 => x"E0823003",
000866 => x"E1510003",
000867 => x"3AFFFFF4",
000868 => x"E2877001",
000869 => x"E5D52030",
000870 => x"E5D53031",
000871 => x"E1833402",
000872 => x"E1570003",
000873 => x"3AFFFFC1",
000874 => x"E3A00000",
000875 => x"E8BD80F0",
000876 => x"00012000",
000877 => x"00012004",
000878 => x"00012020",
000879 => x"E5903000",
000880 => x"E20110FF",
000881 => x"E3530000",
000882 => x"14C31001",
000883 => x"E1A02000",
000884 => x"E1A00001",
000885 => x"15823000",
000886 => x"11A0F00E",
000887 => x"EA00010C",
000888 => x"E92D45F0",
000889 => x"E2525000",
000890 => x"E1A08000",
000891 => x"E1A07001",
000892 => x"C3A02000",
000893 => x"CA000001",
000894 => x"EA000009",
000895 => x"E2822001",
000896 => x"E7D21007",
000897 => x"E3510000",
000898 => x"1AFFFFFB",
000899 => x"E1520005",
000900 => x"A1A05001",
000901 => x"B0625005",
000902 => x"E3130002",
000903 => x"13A0A030",
000904 => x"1A000000",
000905 => x"E3A0A020",
000906 => x"E3130001",
000907 => x"13A06000",
000908 => x"01A04005",
000909 => x"0A000002",
000910 => x"EA00000A",
000911 => x"EBFFFFDE",
000912 => x"E2444001",
000913 => x"E3540000",
000914 => x"E1A00008",
000915 => x"E20A10FF",
000916 => x"CAFFFFF9",
000917 => x"E0646005",
000918 => x"E1A05004",
000919 => x"EA000001",
000920 => x"EBFFFFD5",
000921 => x"E2866001",
000922 => x"E5D73000",
000923 => x"E2531000",
000924 => x"E1A00008",
000925 => x"E2877001",
000926 => x"1AFFFFF8",
000927 => x"EA000001",
000928 => x"EBFFFFCD",
000929 => x"E2866001",
000930 => x"E3550000",
000931 => x"E1A00008",
000932 => x"E20A10FF",
000933 => x"E2455001",
000934 => x"CAFFFFF8",
000935 => x"E1A00006",
000936 => x"E8BD85F0",
000937 => x"E92D4FF0",
000938 => x"E2514000",
000939 => x"E24DD010",
000940 => x"E1A05002",
000941 => x"E1A09000",
000942 => x"E28D6034",
000943 => x"E8960C40",
000944 => x"1A000007",
000945 => x"E3A0C030",
000946 => x"E1A02006",
000947 => x"E1A0300A",
000948 => x"E1A0100D",
000949 => x"E5CDC000",
000950 => x"E5CD4001",
000951 => x"EBFFFFBF",
000952 => x"EA00003C",
000953 => x"E2533000",
000954 => x"13A03001",
000955 => x"E352000A",
000956 => x"13A03000",
000957 => x"E3530000",
000958 => x"0A000003",
000959 => x"E3540000",
000960 => x"B2644000",
000961 => x"B3A08001",
000962 => x"BA000000",
000963 => x"E3A08000",
000964 => x"E3A03000",
000965 => x"E28D700F",
000966 => x"E5CD300F",
000967 => x"EA000010",
000968 => x"E3550010",
000969 => x"0A000002",
000970 => x"EB0000CD",
000971 => x"E0030095",
000972 => x"E0633004",
000973 => x"E3530009",
000974 => x"E083200B",
000975 => x"C242303A",
000976 => x"E2833030",
000977 => x"E3550010",
000978 => x"E1A00004",
000979 => x"E1A01005",
000980 => x"E5673001",
000981 => x"01A04224",
000982 => x"0A000001",
000983 => x"EB0000C0",
000984 => x"E1A04000",
000985 => x"E3540000",
000986 => x"E1A00004",
000987 => x"E1A01005",
000988 => x"E204300F",
000989 => x"1AFFFFE9",
000990 => x"E3580000",
000991 => x"E1A02007",
000992 => x"01A04008",
000993 => x"0A00000D",
000994 => x"E3560000",
000995 => x"0A000007",
000996 => x"E31A0002",
000997 => x"0A000005",
000998 => x"E1A00009",
000999 => x"E3A0102D",
001000 => x"EBFFFF85",
001001 => x"E2466001",
001002 => x"E3A04001",
001003 => x"EA000003",
001004 => x"E3A0302D",
001005 => x"E5423001",
001006 => x"E2477001",
001007 => x"E3A04000",
001008 => x"E1A00009",
001009 => x"E1A01007",
001010 => x"E1A02006",
001011 => x"E1A0300A",
001012 => x"EBFFFF82",
001013 => x"E0840000",
001014 => x"E28DD010",
001015 => x"E8BD8FF0",
001016 => x"E92D41F0",
001017 => x"E1A07000",
001018 => x"E24DD010",
001019 => x"E1A04001",
001020 => x"E1A05002",
001021 => x"E3A06000",
001022 => x"EA00005C",
001023 => x"E3530025",
001024 => x"1A000051",
001025 => x"E5F43001",
001026 => x"E3530000",
001027 => x"0A00005A",
001028 => x"E3530025",
001029 => x"0A000050",
001030 => x"E353002D",
001031 => x"13A08000",
001032 => x"02844001",
001033 => x"03A08001",
001034 => x"EA000001",
001035 => x"E2844001",
001036 => x"E3888002",
001037 => x"E5D43000",
001038 => x"E3530030",
001039 => x"0AFFFFFA",
001040 => x"E3A0E000",
001041 => x"EA000003",
001042 => x"E3A0300A",
001043 => x"E023239E",
001044 => x"E2844001",
001045 => x"E243E030",
001046 => x"E5D42000",
001047 => x"E2423030",
001048 => x"E3530009",
001049 => x"9AFFFFF7",
001050 => x"E3520073",
001051 => x"1A000007",
001052 => x"E4953004",
001053 => x"E59F110C",
001054 => x"E3530000",
001055 => x"11A01003",
001056 => x"E1A0200E",
001057 => x"E1A03008",
001058 => x"E1A00007",
001059 => x"EA00002C",
001060 => x"E3520064",
001061 => x"1A00000A",
001062 => x"E4951004",
001063 => x"E1A00007",
001064 => x"E3A0200A",
001065 => x"E3A03001",
001066 => x"E58DE000",
001067 => x"E58D8004",
001068 => x"E3A0C061",
001069 => x"E58DC008",
001070 => x"EBFFFF79",
001071 => x"E0866000",
001072 => x"EA000029",
001073 => x"E3520078",
001074 => x"04951004",
001075 => x"01A00007",
001076 => x"03A02010",
001077 => x"0A00000E",
001078 => x"E3520058",
001079 => x"1A000007",
001080 => x"E4951004",
001081 => x"E1A00007",
001082 => x"E3A02010",
001083 => x"E3A03000",
001084 => x"E3A0C041",
001085 => x"E58DE000",
001086 => x"E58D8004",
001087 => x"EAFFFFEC",
001088 => x"E3520075",
001089 => x"1A000004",
001090 => x"E4951004",
001091 => x"E1A00007",
001092 => x"E3A0200A",
001093 => x"E3A03000",
001094 => x"EAFFFFE2",
001095 => x"E3520063",
001096 => x"1A000011",
001097 => x"E495C004",
001098 => x"E5CDC00E",
001099 => x"E3A0C000",
001100 => x"E5CDC00F",
001101 => x"E1A0200E",
001102 => x"E1A03008",
001103 => x"E1A00007",
001104 => x"E28D100E",
001105 => x"EBFFFF25",
001106 => x"EAFFFFDB",
001107 => x"E353000A",
001108 => x"01A00007",
001109 => x"03A0100D",
001110 => x"0BFFFF17",
001111 => x"E1A00007",
001112 => x"E5D41000",
001113 => x"EBFFFF14",
001114 => x"E2866001",
001115 => x"E2844001",
001116 => x"E5D43000",
001117 => x"E3530000",
001118 => x"1AFFFF9F",
001119 => x"E1A00006",
001120 => x"E28DD010",
001121 => x"E8BD81F0",
001122 => x"00012058",
001123 => x"E92D000F",
001124 => x"E52DE004",
001125 => x"E24DD004",
001126 => x"E28D0004",
001127 => x"E3A03000",
001128 => x"E5203004",
001129 => x"E59D1008",
001130 => x"E1A0000D",
001131 => x"E28D200C",
001132 => x"EBFFFF8A",
001133 => x"E28DD004",
001134 => x"E49DE004",
001135 => x"E28DD010",
001136 => x"E1A0F00E",
001137 => x"E92D000E",
001138 => x"E52DE004",
001139 => x"E24DD004",
001140 => x"E28D3004",
001141 => x"E5230004",
001142 => x"E59D1008",
001143 => x"E1A0000D",
001144 => x"E28D200C",
001145 => x"EBFFFF7D",
001146 => x"E28DD004",
001147 => x"E49DE004",
001148 => x"E28DD00C",
001149 => x"E1A0F00E",
001150 => x"E59FB46C",
001151 => x"E58B0000",
001152 => x"EAFFFFFC",
001153 => x"E59FB460",
001154 => x"E3A0A011",
001155 => x"E58BA000",
001156 => x"EAFFFFFB",
001157 => x"E59F1454",
001158 => x"E59F3454",
001159 => x"E5932000",
001160 => x"E2022020",
001161 => x"E3520000",
001162 => x"05810000",
001163 => x"01B0F00E",
001164 => x"1AFFFFF9",
001165 => x"E59F2434",
001166 => x"E59F3434",
001167 => x"E1A01580",
001168 => x"E0811480",
001169 => x"E5930000",
001170 => x"E2100010",
001171 => x"05920000",
001172 => x"01A0F00E",
001173 => x"E2511001",
001174 => x"1AFFFFF9",
001175 => x"E3E00000",
001176 => x"E1B0F00E",
001177 => x"E92D4010",
001178 => x"E2002102",
001179 => x"E2013102",
001180 => x"E0224003",
001181 => x"E3100102",
001182 => x"11E00000",
001183 => x"12800001",
001184 => x"E3110102",
001185 => x"11E01001",
001186 => x"12811001",
001187 => x"E1A02001",
001188 => x"E1A01000",
001189 => x"E3520000",
001190 => x"0A000011",
001191 => x"E3A00000",
001192 => x"E3A03001",
001193 => x"E3530000",
001194 => x"03A03201",
001195 => x"0A000003",
001196 => x"E1520001",
001197 => x"91A02082",
001198 => x"91A03083",
001199 => x"9AFFFFF8",
001200 => x"E1510002",
001201 => x"20411002",
001202 => x"20800003",
001203 => x"E1B030A3",
001204 => x"31A020A2",
001205 => x"3AFFFFF9",
001206 => x"E3140102",
001207 => x"11E00000",
001208 => x"12800001",
001209 => x"E8FD8010",
001210 => x"E92D4070",
001211 => x"E1A06000",
001212 => x"E1862001",
001213 => x"E3120003",
001214 => x"1A00002A",
001215 => x"E8B1003C",
001216 => x"E31200FF",
001217 => x"13120CFF",
001218 => x"131208FF",
001219 => x"131204FF",
001220 => x"14862004",
001221 => x"02411004",
001222 => x"131300FF",
001223 => x"13130CFF",
001224 => x"131308FF",
001225 => x"131304FF",
001226 => x"14863004",
001227 => x"02411004",
001228 => x"131400FF",
001229 => x"13140CFF",
001230 => x"131408FF",
001231 => x"131404FF",
001232 => x"14864004",
001233 => x"02411004",
001234 => x"131500FF",
001235 => x"13150CFF",
001236 => x"131508FF",
001237 => x"131504FF",
001238 => x"14865004",
001239 => x"02411004",
001240 => x"1AFFFFE5",
001241 => x"E4913004",
001242 => x"E4C63001",
001243 => x"E21340FF",
001244 => x"08FD8070",
001245 => x"E1A03423",
001246 => x"E4C63001",
001247 => x"E21340FF",
001248 => x"08FD8070",
001249 => x"E1A03423",
001250 => x"E4C63001",
001251 => x"E21340FF",
001252 => x"08FD8070",
001253 => x"E1A03423",
001254 => x"E4C63001",
001255 => x"E21340FF",
001256 => x"08FD8070",
001257 => x"EAFFFFEE",
001258 => x"E4D13001",
001259 => x"E4C63001",
001260 => x"E3530000",
001261 => x"08FD8070",
001262 => x"E4D13001",
001263 => x"E4C63001",
001264 => x"E3530000",
001265 => x"08FD8070",
001266 => x"E4D13001",
001267 => x"E4C63001",
001268 => x"E3530000",
001269 => x"08FD8070",
001270 => x"E4D13001",
001271 => x"E4C63001",
001272 => x"E3530000",
001273 => x"08FD8070",
001274 => x"EAFFFFEE",
001275 => x"E92D41F0",
001276 => x"E1802001",
001277 => x"E3120003",
001278 => x"1A000018",
001279 => x"E8B0001C",
001280 => x"E8B100E0",
001281 => x"E1520005",
001282 => x"1A000012",
001283 => x"01530006",
001284 => x"1A00002B",
001285 => x"01540007",
001286 => x"1A000049",
001287 => x"E31200FF",
001288 => x"13120CFF",
001289 => x"131208FF",
001290 => x"131204FF",
001291 => x"131300FF",
001292 => x"13130CFF",
001293 => x"131308FF",
001294 => x"131304FF",
001295 => x"131400FF",
001296 => x"13140CFF",
001297 => x"131408FF",
001298 => x"131404FF",
001299 => x"1AFFFFEA",
001300 => x"03A00000",
001301 => x"08FD81F0",
001302 => x"E240000C",
001303 => x"E241100C",
001304 => x"E4D02001",
001305 => x"E4D13001",
001306 => x"E0324003",
001307 => x"1A00005A",
001308 => x"E4D05001",
001309 => x"E4D16001",
001310 => x"E3520000",
001311 => x"0A000054",
001312 => x"E0357006",
001313 => x"1A000054",
001314 => x"E4D02001",
001315 => x"E4D13001",
001316 => x"E3550000",
001317 => x"0A00004E",
001318 => x"E0324003",
001319 => x"1A00004E",
001320 => x"E4D05001",
001321 => x"E4D16001",
001322 => x"E3520000",
001323 => x"0A000048",
001324 => x"E0357006",
001325 => x"1A000048",
001326 => x"E3550000",
001327 => x"0A000044",
001328 => x"1AFFFFE6",
001329 => x"E31200FF",
001330 => x"13120CFF",
001331 => x"131208FF",
001332 => x"131204FF",
001333 => x"0A00003E",
001334 => x"E2400008",
001335 => x"E2411008",
001336 => x"E4D02001",
001337 => x"E4D13001",
001338 => x"E0324003",
001339 => x"1A00003A",
001340 => x"E4D05001",
001341 => x"E4D16001",
001342 => x"E3520000",
001343 => x"0A000034",
001344 => x"E0357006",
001345 => x"1A000034",
001346 => x"E4D02001",
001347 => x"E4D13001",
001348 => x"E3550000",
001349 => x"0A00002E",
001350 => x"E0324003",
001351 => x"1A00002E",
001352 => x"E4D05001",
001353 => x"E4D16001",
001354 => x"E3520000",
001355 => x"0A000028",
001356 => x"E0357006",
001357 => x"1A000028",
001358 => x"E3550000",
001359 => x"0A000024",
001360 => x"1AFFFFC6",
001361 => x"E31200FF",
001362 => x"13120CFF",
001363 => x"131208FF",
001364 => x"131204FF",
001365 => x"131300FF",
001366 => x"13130CFF",
001367 => x"131308FF",
001368 => x"131304FF",
001369 => x"0A00001A",
001370 => x"E2400004",
001371 => x"E2411004",
001372 => x"E4D02001",
001373 => x"E4D13001",
001374 => x"E0324003",
001375 => x"1A000016",
001376 => x"E4D05001",
001377 => x"E4D16001",
001378 => x"E3520000",
001379 => x"0A000010",
001380 => x"E0357006",
001381 => x"1A000010",
001382 => x"E4D02001",
001383 => x"E4D13001",
001384 => x"E3550000",
001385 => x"0A00000A",
001386 => x"E0324003",
001387 => x"1A00000A",
001388 => x"E4D05001",
001389 => x"E4D16001",
001390 => x"E3520000",
001391 => x"0A000004",
001392 => x"E0357006",
001393 => x"1A000004",
001394 => x"E3550000",
001395 => x"0A000000",
001396 => x"1AFFFFA2",
001397 => x"03A00000",
001398 => x"08FD81F0",
001399 => x"E0450006",
001400 => x"E8FD81F0",
001401 => x"E59F107C",
001402 => x"E5811000",
001403 => x"E1A0F00E",
001404 => x"E59F1070",
001405 => x"E5910000",
001406 => x"E2800801",
001407 => x"E5810000",
001408 => x"E1A0F00E",
001409 => x"E92D4010",
001410 => x"E3520000",
001411 => x"0A000004",
001412 => x"E0804002",
001413 => x"E4D13001",
001414 => x"E4C03001",
001415 => x"E1500004",
001416 => x"1AFFFFFB",
001417 => x"E8FD8010",
001418 => x"E92D4070",
001419 => x"E3520000",
001420 => x"03A00001",
001421 => x"0A00000A",
001422 => x"E3A03000",
001423 => x"E2833001",
001424 => x"E4D04001",
001425 => x"E4D15001",
001426 => x"E0546005",
001427 => x"11A00006",
001428 => x"1A000003",
001429 => x"E1530002",
001430 => x"03A00000",
001431 => x"0A000000",
001432 => x"EAFFFFF5",
001433 => x"E8FD8070",
001434 => x"07000000",
001435 => x"F0000000",
001436 => x"FFFF0200",
001437 => x"FFFF0218",
001438 => x"E3520007",
001439 => x"E92D45F0",
001440 => x"E1A0C001",
001441 => x"E1A04002",
001442 => x"E1A0A000",
001443 => x"E1A0E000",
001444 => x"83A02000",
001445 => x"8A00001E",
001446 => x"E2443001",
001447 => x"E3530006",
001448 => x"979FF103",
001449 => x"EA000140",
001450 => x"000116FC",
001451 => x"000116F4",
001452 => x"000116EC",
001453 => x"000116E4",
001454 => x"000116DC",
001455 => x"000116D4",
001456 => x"000116C4",
001457 => x"E4D13001",
001458 => x"E1A0E000",
001459 => x"E4CE3001",
001460 => x"E1A0C001",
001461 => x"E4DC3001",
001462 => x"E4CE3001",
001463 => x"E4DC3001",
001464 => x"E4CE3001",
001465 => x"E4DC3001",
001466 => x"E4CE3001",
001467 => x"E4DC3001",
001468 => x"E4CE3001",
001469 => x"E4DC3001",
001470 => x"E4CE3001",
001471 => x"E5DC3000",
001472 => x"E5CE3000",
001473 => x"EA000128",
001474 => x"E7D23001",
001475 => x"E7C2300A",
001476 => x"E2822001",
001477 => x"E08AE002",
001478 => x"E31E0003",
001479 => x"1AFFFFF9",
001480 => x"E0811002",
001481 => x"E2013003",
001482 => x"E0626004",
001483 => x"E3530003",
001484 => x"979FF103",
001485 => x"EA00011B",
001486 => x"00011748",
001487 => x"00011818",
001488 => x"00011928",
001489 => x"00011A38",
001490 => x"E1A02126",
001491 => x"E3A0C000",
001492 => x"EA000003",
001493 => x"E79C3001",
001494 => x"E2422001",
001495 => x"E78C300E",
001496 => x"E28CC004",
001497 => x"E3120007",
001498 => x"1AFFFFF9",
001499 => x"E08E500C",
001500 => x"E081100C",
001501 => x"E1A021A2",
001502 => x"E1A0E005",
001503 => x"E1A0C001",
001504 => x"E1A04002",
001505 => x"EA00000F",
001506 => x"E51C3020",
001507 => x"E50E3020",
001508 => x"E51C301C",
001509 => x"E50E301C",
001510 => x"E51C3018",
001511 => x"E50E3018",
001512 => x"E51C3014",
001513 => x"E50E3014",
001514 => x"E51C3010",
001515 => x"E50E3010",
001516 => x"E51C300C",
001517 => x"E50E300C",
001518 => x"E51C3008",
001519 => x"E50E3008",
001520 => x"E51C3004",
001521 => x"E50E3004",
001522 => x"E2444001",
001523 => x"E3740001",
001524 => x"E28EE020",
001525 => x"E28CC020",
001526 => x"1AFFFFEA",
001527 => x"E2063003",
001528 => x"E1A02282",
001529 => x"E2433001",
001530 => x"E085C002",
001531 => x"E0811002",
001532 => x"E3530006",
001533 => x"979FF103",
001534 => x"EA0000EB",
001535 => x"00011B9C",
001536 => x"00011B94",
001537 => x"00011B8C",
001538 => x"00011B84",
001539 => x"00011B7C",
001540 => x"00011B74",
001541 => x"00011B6C",
001542 => x"E3C10003",
001543 => x"E5904000",
001544 => x"E3CE1003",
001545 => x"E1A0C126",
001546 => x"E1A02001",
001547 => x"EA000003",
001548 => x"E7954003",
001549 => x"E18E3C04",
001550 => x"E5023004",
001551 => x"E24CC001",
001552 => x"E2822004",
001553 => x"E31C0007",
001554 => x"E2615000",
001555 => x"E1A0E424",
001556 => x"E0803002",
001557 => x"1AFFFFF5",
001558 => x"E0613000",
001559 => x"E0837002",
001560 => x"E1A001AC",
001561 => x"E2428004",
001562 => x"E1A0E008",
001563 => x"E1A0C007",
001564 => x"E1A05000",
001565 => x"EA00001F",
001566 => x"E51C2020",
001567 => x"E1A03C02",
001568 => x"E1833424",
001569 => x"E50E3020",
001570 => x"E51C101C",
001571 => x"E1A03C01",
001572 => x"E1833422",
001573 => x"E50E301C",
001574 => x"E51C2018",
001575 => x"E1A03C02",
001576 => x"E1833421",
001577 => x"E50E3018",
001578 => x"E51C1014",
001579 => x"E1A03C01",
001580 => x"E1833422",
001581 => x"E50E3014",
001582 => x"E51C2010",
001583 => x"E1A03C02",
001584 => x"E1833421",
001585 => x"E50E3010",
001586 => x"E51C100C",
001587 => x"E1A03C01",
001588 => x"E1833422",
001589 => x"E50E300C",
001590 => x"E51C2008",
001591 => x"E1A03C02",
001592 => x"E1833421",
001593 => x"E50E3008",
001594 => x"E51C4004",
001595 => x"E1A03C04",
001596 => x"E1833422",
001597 => x"E50E3004",
001598 => x"E2455001",
001599 => x"E3750001",
001600 => x"E28EE020",
001601 => x"E28CC020",
001602 => x"1AFFFFDA",
001603 => x"E1A03280",
001604 => x"E2062003",
001605 => x"E0871003",
001606 => x"E2422001",
001607 => x"E088C003",
001608 => x"E2411003",
001609 => x"EA000086",
001610 => x"E3C10003",
001611 => x"E5904000",
001612 => x"E3CE1003",
001613 => x"E1A0C126",
001614 => x"E1A02001",
001615 => x"EA000003",
001616 => x"E7954003",
001617 => x"E18E3804",
001618 => x"E5023004",
001619 => x"E24CC001",
001620 => x"E2822004",
001621 => x"E31C0007",
001622 => x"E2615000",
001623 => x"E1A0E824",
001624 => x"E0803002",
001625 => x"1AFFFFF5",
001626 => x"E0613000",
001627 => x"E0837002",
001628 => x"E1A001AC",
001629 => x"E2428004",
001630 => x"E1A0E008",
001631 => x"E1A0C007",
001632 => x"E1A05000",
001633 => x"EA00001F",
001634 => x"E51C2020",
001635 => x"E1A03802",
001636 => x"E1833824",
001637 => x"E50E3020",
001638 => x"E51C101C",
001639 => x"E1A03801",
001640 => x"E1833822",
001641 => x"E50E301C",
001642 => x"E51C2018",
001643 => x"E1A03802",
001644 => x"E1833821",
001645 => x"E50E3018",
001646 => x"E51C1014",
001647 => x"E1A03801",
001648 => x"E1833822",
001649 => x"E50E3014",
001650 => x"E51C2010",
001651 => x"E1A03802",
001652 => x"E1833821",
001653 => x"E50E3010",
001654 => x"E51C100C",
001655 => x"E1A03801",
001656 => x"E1833822",
001657 => x"E50E300C",
001658 => x"E51C2008",
001659 => x"E1A03802",
001660 => x"E1833821",
001661 => x"E50E3008",
001662 => x"E51C4004",
001663 => x"E1A03804",
001664 => x"E1833822",
001665 => x"E50E3004",
001666 => x"E2455001",
001667 => x"E3750001",
001668 => x"E28EE020",
001669 => x"E28CC020",
001670 => x"1AFFFFDA",
001671 => x"E1A03280",
001672 => x"E2062003",
001673 => x"E0871003",
001674 => x"E2422001",
001675 => x"E088C003",
001676 => x"E2411002",
001677 => x"EA000042",
001678 => x"E3C10003",
001679 => x"E5904000",
001680 => x"E3CE1003",
001681 => x"E1A0C126",
001682 => x"E1A02001",
001683 => x"EA000003",
001684 => x"E7954003",
001685 => x"E18E3404",
001686 => x"E5023004",
001687 => x"E24CC001",
001688 => x"E2822004",
001689 => x"E31C0007",
001690 => x"E2615000",
001691 => x"E1A0EC24",
001692 => x"E0803002",
001693 => x"1AFFFFF5",
001694 => x"E0613000",
001695 => x"E0837002",
001696 => x"E1A001AC",
001697 => x"E2428004",
001698 => x"E1A0E008",
001699 => x"E1A0C007",
001700 => x"E1A05000",
001701 => x"EA00001F",
001702 => x"E51C2020",
001703 => x"E1A03402",
001704 => x"E1833C24",
001705 => x"E50E3020",
001706 => x"E51C101C",
001707 => x"E1A03401",
001708 => x"E1833C22",
001709 => x"E50E301C",
001710 => x"E51C2018",
001711 => x"E1A03402",
001712 => x"E1833C21",
001713 => x"E50E3018",
001714 => x"E51C1014",
001715 => x"E1A03401",
001716 => x"E1833C22",
001717 => x"E50E3014",
001718 => x"E51C2010",
001719 => x"E1A03402",
001720 => x"E1833C21",
001721 => x"E50E3010",
001722 => x"E51C100C",
001723 => x"E1A03401",
001724 => x"E1833C22",
001725 => x"E50E300C",
001726 => x"E51C2008",
001727 => x"E1A03402",
001728 => x"E1833C21",
001729 => x"E50E3008",
001730 => x"E51C4004",
001731 => x"E1A03404",
001732 => x"E1833C22",
001733 => x"E50E3004",
001734 => x"E2455001",
001735 => x"E3750001",
001736 => x"E28EE020",
001737 => x"E28CC020",
001738 => x"1AFFFFDA",
001739 => x"E1A03280",
001740 => x"E2062003",
001741 => x"E0871003",
001742 => x"E2422001",
001743 => x"E088C003",
001744 => x"E2411001",
001745 => x"E3520006",
001746 => x"979FF102",
001747 => x"EA000016",
001748 => x"00011B9C",
001749 => x"00011B94",
001750 => x"00011B8C",
001751 => x"00011B84",
001752 => x"00011B7C",
001753 => x"00011B74",
001754 => x"00011B6C",
001755 => x"E4D13001",
001756 => x"E4CC3001",
001757 => x"E4D13001",
001758 => x"E4CC3001",
001759 => x"E4D13001",
001760 => x"E4CC3001",
001761 => x"E4D13001",
001762 => x"E4CC3001",
001763 => x"E4D13001",
001764 => x"E4CC3001",
001765 => x"E4D13001",
001766 => x"E4CC3001",
001767 => x"E5D13000",
001768 => x"E5CC3000",
001769 => x"EA000000",
001770 => x"E8BD85F0",
001771 => x"E1A0000A",
001772 => x"E8BD85F0",
001773 => x"00001021",
001774 => x"20423063",
001775 => x"408450A5",
001776 => x"60C670E7",
001777 => x"81089129",
001778 => x"A14AB16B",
001779 => x"C18CD1AD",
001780 => x"E1CEF1EF",
001781 => x"12310210",
001782 => x"32732252",
001783 => x"52B54294",
001784 => x"72F762D6",
001785 => x"93398318",
001786 => x"B37BA35A",
001787 => x"D3BDC39C",
001788 => x"F3FFE3DE",
001789 => x"24623443",
001790 => x"04201401",
001791 => x"64E674C7",
001792 => x"44A45485",
001793 => x"A56AB54B",
001794 => x"85289509",
001795 => x"E5EEF5CF",
001796 => x"C5ACD58D",
001797 => x"36532672",
001798 => x"16110630",
001799 => x"76D766F6",
001800 => x"569546B4",
001801 => x"B75BA77A",
001802 => x"97198738",
001803 => x"F7DFE7FE",
001804 => x"D79DC7BC",
001805 => x"48C458E5",
001806 => x"688678A7",
001807 => x"08401861",
001808 => x"28023823",
001809 => x"C9CCD9ED",
001810 => x"E98EF9AF",
001811 => x"89489969",
001812 => x"A90AB92B",
001813 => x"5AF54AD4",
001814 => x"7AB76A96",
001815 => x"1A710A50",
001816 => x"3A332A12",
001817 => x"DBFDCBDC",
001818 => x"FBBFEB9E",
001819 => x"9B798B58",
001820 => x"BB3BAB1A",
001821 => x"6CA67C87",
001822 => x"4CE45CC5",
001823 => x"2C223C03",
001824 => x"0C601C41",
001825 => x"EDAEFD8F",
001826 => x"CDECDDCD",
001827 => x"AD2ABD0B",
001828 => x"8D689D49",
001829 => x"7E976EB6",
001830 => x"5ED54EF4",
001831 => x"3E132E32",
001832 => x"1E510E70",
001833 => x"FF9FEFBE",
001834 => x"DFDDCFFC",
001835 => x"BF1BAF3A",
001836 => x"9F598F78",
001837 => x"918881A9",
001838 => x"B1CAA1EB",
001839 => x"D10CC12D",
001840 => x"F14EE16F",
001841 => x"108000A1",
001842 => x"30C220E3",
001843 => x"50044025",
001844 => x"70466067",
001845 => x"83B99398",
001846 => x"A3FBB3DA",
001847 => x"C33DD31C",
001848 => x"E37FF35E",
001849 => x"02B11290",
001850 => x"22F332D2",
001851 => x"42355214",
001852 => x"62777256",
001853 => x"B5EAA5CB",
001854 => x"95A88589",
001855 => x"F56EE54F",
001856 => x"D52CC50D",
001857 => x"34E224C3",
001858 => x"14A00481",
001859 => x"74666447",
001860 => x"54244405",
001861 => x"A7DBB7FA",
001862 => x"879997B8",
001863 => x"E75FF77E",
001864 => x"C71DD73C",
001865 => x"26D336F2",
001866 => x"069116B0",
001867 => x"66577676",
001868 => x"46155634",
001869 => x"D94CC96D",
001870 => x"F90EE92F",
001871 => x"99C889E9",
001872 => x"B98AA9AB",
001873 => x"58444865",
001874 => x"78066827",
001875 => x"18C008E1",
001876 => x"388228A3",
001877 => x"CB7DDB5C",
001878 => x"EB3FFB1E",
001879 => x"8BF99BD8",
001880 => x"ABBBBB9A",
001881 => x"4A755A54",
001882 => x"6A377A16",
001883 => x"0AF11AD0",
001884 => x"2AB33A92",
001885 => x"FD2EED0F",
001886 => x"DD6CCD4D",
001887 => x"BDAAAD8B",
001888 => x"9DE88DC9",
001889 => x"7C266C07",
001890 => x"5C644C45",
001891 => x"3CA22C83",
001892 => x"1CE00CC1",
001893 => x"EF1FFF3E",
001894 => x"CF5DDF7C",
001895 => x"AF9BBFBA",
001896 => x"8FD99FF8",
001897 => x"6E177E36",
001898 => x"4E555E74",
001899 => x"2E933EB2",
001900 => x"0ED11EF0",
001901 => x"20000000",
001902 => x"436F6D6D",
001903 => x"616E6473",
001904 => x"0A000000",
001905 => x"6C000000",
001906 => x"3A204C6F",
001907 => x"61642065",
001908 => x"6C662066",
001909 => x"696C650A",
001910 => x"00000000",
001911 => x"62203C61",
001912 => x"64647265",
001913 => x"73733E00",
001914 => x"3A204C6F",
001915 => x"61642062",
001916 => x"696E6172",
001917 => x"79206669",
001918 => x"6C652074",
001919 => x"6F203C61",
001920 => x"64647265",
001921 => x"73733E0A",
001922 => x"00000000",
001923 => x"64203C73",
001924 => x"74617274",
001925 => x"20616464",
001926 => x"72657373",
001927 => x"3E203C6E",
001928 => x"756D2062",
001929 => x"79746573",
001930 => x"3E203A20",
001931 => x"44756D70",
001932 => x"206D656D",
001933 => x"0A000000",
001934 => x"68000000",
001935 => x"3A205072",
001936 => x"696E7420",
001937 => x"68656C70",
001938 => x"206D6573",
001939 => x"73616765",
001940 => x"0A000000",
001941 => x"6A203C61",
001942 => x"64647265",
001943 => x"73733E00",
001944 => x"3A204578",
001945 => x"65637574",
001946 => x"65206C6F",
001947 => x"61646564",
001948 => x"20656C66",
001949 => x"2C206A75",
001950 => x"6D70696E",
001951 => x"6720746F",
001952 => x"203C6164",
001953 => x"64726573",
001954 => x"733E0A00",
001955 => x"70203C61",
001956 => x"64647265",
001957 => x"73733E00",
001958 => x"3A205072",
001959 => x"696E7420",
001960 => x"61736369",
001961 => x"69206D65",
001962 => x"6D20756E",
001963 => x"74696C20",
001964 => x"66697273",
001965 => x"7420300A",
001966 => x"00000000",
001967 => x"72203C61",
001968 => x"64647265",
001969 => x"73733E00",
001970 => x"3A205265",
001971 => x"6164206D",
001972 => x"656D0A00",
001973 => x"73000000",
001974 => x"3A20436F",
001975 => x"72652073",
001976 => x"74617475",
001977 => x"730A0000",
001978 => x"77203C61",
001979 => x"64647265",
001980 => x"73733E20",
001981 => x"3C76616C",
001982 => x"75653E00",
001983 => x"3A205772",
001984 => x"69746520",
001985 => x"6D656D0A",
001986 => x"00000000",
001987 => x"6D656D20",
001988 => x"30782530",
001989 => x"3878203D",
001990 => x"20307825",
001991 => x"3038780A",
001992 => x"00000000",
001993 => x"25730A00",
001994 => x"53656E64",
001995 => x"2066696C",
001996 => x"6520772F",
001997 => x"20314B20",
001998 => x"586D6F64",
001999 => x"656D2070",
002000 => x"726F746F",
002001 => x"636F6C20",
002002 => x"66726F6D",
002003 => x"20746572",
002004 => x"6D696E61",
002005 => x"6C20656D",
002006 => x"756C6174",
002007 => x"6F72206E",
002008 => x"6F772E2E",
002009 => x"2E000000",
002010 => x"586D6F64",
002011 => x"656D2065",
002012 => x"72726F72",
002013 => x"2066696C",
002014 => x"65207369",
002015 => x"7A652030",
002016 => x"78257820",
002017 => x"0A000000",
002018 => x"0A656C66",
002019 => x"2073706C",
002020 => x"69740A00",
002021 => x"6A203078",
002022 => x"25303878",
002023 => x"0A000000",
002024 => x"496E7661",
002025 => x"6C696420",
002026 => x"636F6D6D",
002027 => x"616E6400",
002028 => x"2563416D",
002029 => x"62657220",
002030 => x"426F6F74",
002031 => x"204C6F61",
002032 => x"64657220",
002033 => x"77697468",
002034 => x"20444530",
002035 => x"2D4E414E",
002036 => x"4F203332",
002037 => x"4D422073",
002038 => x"7570706F",
002039 => x"72747625",
002040 => x"730A0000",
002041 => x"32303135",
002042 => x"2D31302D",
002043 => x"30330000",
002044 => x"52656164",
002045 => x"790A3E20",
002046 => x"00000000",
002047 => x"3E200000",
002048 => x"454C4600",
002049 => x"4552524F",
002050 => x"523A204E",
002051 => x"6F742061",
002052 => x"6E20454C",
002053 => x"46206669",
002054 => x"6C652E0A",
002055 => x"00000000",
002056 => x"4552524F",
002057 => x"523A2045",
002058 => x"4C462066",
002059 => x"696C6520",
002060 => x"6E6F7420",
002061 => x"74617267",
002062 => x"65747469",
002063 => x"6E672063",
002064 => x"6F727265",
002065 => x"63742070",
002066 => x"726F6365",
002067 => x"73736F72",
002068 => x"20747970",
002069 => x"650A0000",
002070 => x"286E756C",
002071 => x"6C290000",
others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;